module mux_8 ( ctrl0, ctrl1, ctrl2, ctrl3, ctrl4, ctrl5, ctrl6, ctrl7, in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, in64, in65, in66, in67, in68, in69, in70, in71, in72, in73, in74, in75, in76, in77, in78, in79, in80, in81, in82, in83, in84, in85, in86, in87, in88, in89, in90, in91, in92, in93, in94, in95, in96, in97, in98, in99, in100, in101, in102, in103, in104, in105, in106, in107, in108, in109, in110, in111, in112, in113, in114, in115, in116, in117, in118, in119, in120, in121, in122, in123, in124, in125, in126, in127, in128, in129, in130, in131, in132, in133, in134, in135, in136, in137, in138, in139, in140, in141, in142, in143, in144, in145, in146, in147, in148, in149, in150, in151, in152, in153, in154, in155, in156, in157, in158, in159, in160, in161, in162, in163, in164, in165, in166, in167, in168, in169, in170, in171, in172, in173, in174, in175, in176, in177, in178, in179, in180, in181, in182, in183, in184, in185, in186, in187, in188, in189, in190, in191, in192, in193, in194, in195, in196, in197, in198, in199, in200, in201, in202, in203, in204, in205, in206, in207, in208, in209, in210, in211, in212, in213, in214, in215, in216, in217, in218, in219, in220, in221, in222, in223, in224, in225, in226, in227, in228, in229, in230, in231, in232, in233, in234, in235, in236, in237, in238, in239, in240, in241, in242, in243, in244, in245, in246, in247, in248, in249, in250, in251, in252, in253, in254, in255, out);
input ctrl0, ctrl1, ctrl2, ctrl3, ctrl4, ctrl5, ctrl6, ctrl7, in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, in64, in65, in66, in67, in68, in69, in70, in71, in72, in73, in74, in75, in76, in77, in78, in79, in80, in81, in82, in83, in84, in85, in86, in87, in88, in89, in90, in91, in92, in93, in94, in95, in96, in97, in98, in99, in100, in101, in102, in103, in104, in105, in106, in107, in108, in109, in110, in111, in112, in113, in114, in115, in116, in117, in118, in119, in120, in121, in122, in123, in124, in125, in126, in127, in128, in129, in130, in131, in132, in133, in134, in135, in136, in137, in138, in139, in140, in141, in142, in143, in144, in145, in146, in147, in148, in149, in150, in151, in152, in153, in154, in155, in156, in157, in158, in159, in160, in161, in162, in163, in164, in165, in166, in167, in168, in169, in170, in171, in172, in173, in174, in175, in176, in177, in178, in179, in180, in181, in182, in183, in184, in185, in186, in187, in188, in189, in190, in191, in192, in193, in194, in195, in196, in197, in198, in199, in200, in201, in202, in203, in204, in205, in206, in207, in208, in209, in210, in211, in212, in213, in214, in215, in216, in217, in218, in219, in220, in221, in222, in223, in224, in225, in226, in227, in228, in229, in230, in231, in232, in233, in234, in235, in236, in237, in238, in239, in240, in241, in242, in243, in244, in245, in246, in247, in248, in249, in250, in251, in252, in253, in254, in255;
output out;
assign out = ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7  ) ? in1 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7  ) ? in2 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7  ) ? in3 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7  ) ? in4 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7  ) ? in5 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7  ) ? in6 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7  ) ? in7 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7  ) ? in8 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7  ) ? in9 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7  ) ? in10 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7  ) ? in11 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7  ) ? in12 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7  ) ? in13 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7  ) ? in14 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7  ) ? in15 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7  ) ? in16 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7  ) ? in17 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7  ) ? in18 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7  ) ? in19 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7  ) ? in20 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7  ) ? in21 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7  ) ? in22 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7  ) ? in23 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7  ) ? in24 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7  ) ? in25 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7  ) ? in26 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7  ) ? in27 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7  ) ? in28 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7  ) ? in29 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7  ) ? in30 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7  ) ? in31 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7  ) ? in32 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7  ) ? in33 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7  ) ? in34 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7  ) ? in35 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7  ) ? in36 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7  ) ? in37 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7  ) ? in38 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7  ) ? in39 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7  ) ? in40 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7  ) ? in41 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7  ) ? in42 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7  ) ? in43 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7  ) ? in44 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7  ) ? in45 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7  ) ? in46 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7  ) ? in47 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7  ) ? in48 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7  ) ? in49 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7  ) ? in50 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7  ) ? in51 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7  ) ? in52 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7  ) ? in53 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7  ) ? in54 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7  ) ? in55 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7  ) ? in56 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7  ) ? in57 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7  ) ? in58 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7  ) ? in59 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7  ) ? in60 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7  ) ? in61 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7  ) ? in62 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7  ) ? in63 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7  ) ? in64 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7  ) ? in65 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7  ) ? in66 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7  ) ? in67 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7  ) ? in68 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7  ) ? in69 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7  ) ? in70 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7  ) ? in71 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7  ) ? in72 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7  ) ? in73 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7  ) ? in74 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7  ) ? in75 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7  ) ? in76 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7  ) ? in77 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7  ) ? in78 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7  ) ? in79 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7  ) ? in80 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7  ) ? in81 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7  ) ? in82 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7  ) ? in83 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7  ) ? in84 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7  ) ? in85 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7  ) ? in86 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7  ) ? in87 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7  ) ? in88 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7  ) ? in89 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7  ) ? in90 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7  ) ? in91 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7  ) ? in92 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7  ) ? in93 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7  ) ? in94 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7  ) ? in95 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7  ) ? in96 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7  ) ? in97 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7  ) ? in98 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7  ) ? in99 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7  ) ? in100 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7  ) ? in101 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7  ) ? in102 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7  ) ? in103 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7  ) ? in104 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7  ) ? in105 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7  ) ? in106 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7  ) ? in107 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7  ) ? in108 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7  ) ? in109 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7  ) ? in110 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7  ) ? in111 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7  ) ? in112 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7  ) ? in113 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7  ) ? in114 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7  ) ? in115 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7  ) ? in116 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7  ) ? in117 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7  ) ? in118 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7  ) ? in119 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7  ) ? in120 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7  ) ? in121 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7  ) ? in122 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7  ) ? in123 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7  ) ? in124 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7  ) ? in125 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7  ) ? in126 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7  ) ? in127 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7  ) ? in128 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7  ) ? in129 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7  ) ? in130 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7  ) ? in131 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7  ) ? in132 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7  ) ? in133 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7  ) ? in134 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7  ) ? in135 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7  ) ? in136 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7  ) ? in137 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7  ) ? in138 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7  ) ? in139 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7  ) ? in140 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7  ) ? in141 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7  ) ? in142 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7  ) ? in143 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7  ) ? in144 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7  ) ? in145 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7  ) ? in146 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7  ) ? in147 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7  ) ? in148 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7  ) ? in149 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7  ) ? in150 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7  ) ? in151 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7  ) ? in152 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7  ) ? in153 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7  ) ? in154 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7  ) ? in155 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7  ) ? in156 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7  ) ? in157 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7  ) ? in158 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7  ) ? in159 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7  ) ? in160 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7  ) ? in161 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7  ) ? in162 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7  ) ? in163 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7  ) ? in164 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7  ) ? in165 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7  ) ? in166 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7  ) ? in167 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7  ) ? in168 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7  ) ? in169 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7  ) ? in170 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7  ) ? in171 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7  ) ? in172 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7  ) ? in173 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7  ) ? in174 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7  ) ? in175 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7  ) ? in176 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7  ) ? in177 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7  ) ? in178 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7  ) ? in179 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7  ) ? in180 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7  ) ? in181 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7  ) ? in182 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7  ) ? in183 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7  ) ? in184 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7  ) ? in185 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7  ) ? in186 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7  ) ? in187 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7  ) ? in188 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7  ) ? in189 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7  ) ? in190 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7  ) ? in191 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7  ) ? in192 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7  ) ? in193 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7  ) ? in194 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7  ) ? in195 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7  ) ? in196 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7  ) ? in197 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7  ) ? in198 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7  ) ? in199 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7  ) ? in200 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7  ) ? in201 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7  ) ? in202 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7  ) ? in203 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7  ) ? in204 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7  ) ? in205 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7  ) ? in206 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7  ) ? in207 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7  ) ? in208 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7  ) ? in209 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7  ) ? in210 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7  ) ? in211 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7  ) ? in212 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7  ) ? in213 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7  ) ? in214 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7  ) ? in215 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7  ) ? in216 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7  ) ? in217 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7  ) ? in218 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7  ) ? in219 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7  ) ? in220 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7  ) ? in221 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7  ) ? in222 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7  ) ? in223 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7  ) ? in224 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7  ) ? in225 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7  ) ? in226 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7  ) ? in227 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7  ) ? in228 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7  ) ? in229 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7  ) ? in230 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7  ) ? in231 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7  ) ? in232 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7  ) ? in233 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7  ) ? in234 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7  ) ? in235 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7  ) ? in236 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7  ) ? in237 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7  ) ? in238 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7  ) ? in239 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7  ) ? in240 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7  ) ? in241 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7  ) ? in242 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7  ) ? in243 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7  ) ? in244 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7  ) ? in245 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7  ) ? in246 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7  ) ? in247 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7  ) ? in248 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7  ) ? in249 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7  ) ? in250 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7  ) ? in251 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7  ) ? in252 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7  ) ? in253 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7  ) ? in254 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7  ) ? in255 : 
             in0;
endmodule
