module mux_7 ( ctrl0, ctrl1, ctrl2, ctrl3, ctrl4, ctrl5, ctrl6, in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, in64, in65, in66, in67, in68, in69, in70, in71, in72, in73, in74, in75, in76, in77, in78, in79, in80, in81, in82, in83, in84, in85, in86, in87, in88, in89, in90, in91, in92, in93, in94, in95, in96, in97, in98, in99, in100, in101, in102, in103, in104, in105, in106, in107, in108, in109, in110, in111, in112, in113, in114, in115, in116, in117, in118, in119, in120, in121, in122, in123, in124, in125, in126, in127, out);
input ctrl0, ctrl1, ctrl2, ctrl3, ctrl4, ctrl5, ctrl6, in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, in64, in65, in66, in67, in68, in69, in70, in71, in72, in73, in74, in75, in76, in77, in78, in79, in80, in81, in82, in83, in84, in85, in86, in87, in88, in89, in90, in91, in92, in93, in94, in95, in96, in97, in98, in99, in100, in101, in102, in103, in104, in105, in106, in107, in108, in109, in110, in111, in112, in113, in114, in115, in116, in117, in118, in119, in120, in121, in122, in123, in124, in125, in126, in127;
output out;
assign out = ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6  ) ? in1 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6  ) ? in2 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6  ) ? in3 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6  ) ? in4 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6  ) ? in5 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6  ) ? in6 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6  ) ? in7 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6  ) ? in8 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6  ) ? in9 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6  ) ? in10 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6  ) ? in11 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6  ) ? in12 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6  ) ? in13 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6  ) ? in14 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6  ) ? in15 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6  ) ? in16 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6  ) ? in17 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6  ) ? in18 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6  ) ? in19 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6  ) ? in20 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6  ) ? in21 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6  ) ? in22 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6  ) ? in23 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6  ) ? in24 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6  ) ? in25 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6  ) ? in26 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6  ) ? in27 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6  ) ? in28 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6  ) ? in29 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6  ) ? in30 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6  ) ? in31 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6  ) ? in32 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6  ) ? in33 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6  ) ? in34 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6  ) ? in35 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6  ) ? in36 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6  ) ? in37 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6  ) ? in38 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6  ) ? in39 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6  ) ? in40 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6  ) ? in41 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6  ) ? in42 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6  ) ? in43 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6  ) ? in44 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6  ) ? in45 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6  ) ? in46 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6  ) ? in47 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6  ) ? in48 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6  ) ? in49 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6  ) ? in50 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6  ) ? in51 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6  ) ? in52 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6  ) ? in53 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6  ) ? in54 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6  ) ? in55 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6  ) ? in56 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6  ) ? in57 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6  ) ? in58 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6  ) ? in59 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6  ) ? in60 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6  ) ? in61 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6  ) ? in62 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6  ) ? in63 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6  ) ? in64 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6  ) ? in65 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6  ) ? in66 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6  ) ? in67 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6  ) ? in68 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6  ) ? in69 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6  ) ? in70 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6  ) ? in71 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6  ) ? in72 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6  ) ? in73 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6  ) ? in74 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6  ) ? in75 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6  ) ? in76 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6  ) ? in77 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6  ) ? in78 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6  ) ? in79 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6  ) ? in80 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6  ) ? in81 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6  ) ? in82 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6  ) ? in83 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6  ) ? in84 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6  ) ? in85 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6  ) ? in86 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6  ) ? in87 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6  ) ? in88 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6  ) ? in89 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6  ) ? in90 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6  ) ? in91 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6  ) ? in92 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6  ) ? in93 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6  ) ? in94 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6  ) ? in95 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6  ) ? in96 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6  ) ? in97 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6  ) ? in98 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6  ) ? in99 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6  ) ? in100 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6  ) ? in101 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6  ) ? in102 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6  ) ? in103 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6  ) ? in104 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6  ) ? in105 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6  ) ? in106 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6  ) ? in107 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6  ) ? in108 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6  ) ? in109 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6  ) ? in110 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6  ) ? in111 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6  ) ? in112 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6  ) ? in113 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6  ) ? in114 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6  ) ? in115 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6  ) ? in116 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6  ) ? in117 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6  ) ? in118 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6  ) ? in119 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6  ) ? in120 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6  ) ? in121 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6  ) ? in122 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6  ) ? in123 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6  ) ? in124 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6  ) ? in125 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6  ) ? in126 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6  ) ? in127 : 
             in0;
endmodule
