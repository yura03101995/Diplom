// Benchmark "top" written by ABC on Mon Apr 24 11:13:58 2017

module top ( 
    in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13,
    in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25,
    in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37,
    in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49,
    in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61,
    in62, in63, in64, in65, in66, in67, in68, in69, in70, in71, in72, in73,
    in74, in75, in76, in77, in78, in79, in80, in81, in82, in83, in84, in85,
    in86, in87, in88, in89, in90, in91, in92, in93, in94, in95, in96, in97,
    in98, in99, in100, in101, in102, in103, in104, in105, in106, in107,
    in108, in109, in110, in111, in112, in113, in114,
    out1  );
  input  in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12,
    in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24,
    in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36,
    in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48,
    in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60,
    in61, in62, in63, in64, in65, in66, in67, in68, in69, in70, in71, in72,
    in73, in74, in75, in76, in77, in78, in79, in80, in81, in82, in83, in84,
    in85, in86, in87, in88, in89, in90, in91, in92, in93, in94, in95, in96,
    in97, in98, in99, in100, in101, in102, in103, in104, in105, in106,
    in107, in108, in109, in110, in111, in112, in113, in114;
  output out1;
  wire n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
    n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
    n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
    n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
    n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
    n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
    n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
    n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
    n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
    n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
    n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
    n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
    n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
    n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
    n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
    n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
    n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
    n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
    n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
    n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
    n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
    n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
    n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
    n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
    n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
    n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
    n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
    n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
    n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
    n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
    n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
    n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
    n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
    n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
    n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
    n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
    n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
    n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
    n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
    n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
    n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
    n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
    n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
    n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
    n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
    n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
    n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
    n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
    n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
    n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
    n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
    n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
    n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
    n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
    n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
    n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
    n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
    n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
    n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
    n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
    n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
    n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
    n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
    n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
    n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
    n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
    n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
    n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
    n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
    n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
    n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
    n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
    n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
    n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
    n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
    n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
    n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
    n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
    n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
    n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
    n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
    n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
    n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
    n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
    n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
    n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
    n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
    n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
    n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
    n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
    n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
    n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
    n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
    n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
    n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
    n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
    n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
    n1262;
  not    g0000(.a(in7), .O(n116));
  not    g0001(.a(in75), .O(n117));
  xnor2a g0002(.a(in97), .b(in14), .O(n118));
  nand3  g0003(.a(in83), .b(in55), .c(in35), .O(n119));
  nand3  g0004(.a(n119), .b(n118), .c(in40), .O(n120));
  nand2  g0005(.a(n120), .b(n117), .O(n121));
  xor2a  g0006(.a(n121), .b(n116), .O(n122));
  not    g0007(.a(in101), .O(n123));
  not    g0008(.a(in54), .O(n124));
  not    g0009(.a(in93), .O(n125));
  nand3  g0010(.a(in112), .b(n125), .c(n124), .O(n126));
  nand3  g0011(.a(in83), .b(in10), .c(in2), .O(n127));
  xor2a  g0012(.a(in106), .b(in41), .O(n128));
  xor2a  g0013(.a(n128), .b(n127), .O(n129));
  nand3  g0014(.a(n129), .b(n126), .c(in64), .O(n130));
  not    g0015(.a(in71), .O(n131));
  not    g0016(.a(in31), .O(n132));
  not    g0017(.a(in42), .O(n133));
  nand4  g0018(.a(in65), .b(in45), .c(n133), .d(n132), .O(n134));
  nand3  g0019(.a(n134), .b(n131), .c(in51), .O(n135));
  nand3  g0020(.a(n135), .b(n130), .c(in65), .O(n136));
  not    g0021(.a(in5), .O(n137));
  not    g0022(.a(in1), .O(n138));
  not    g0023(.a(in58), .O(n139));
  not    g0024(.a(in111), .O(n140));
  nand3  g0025(.a(n140), .b(n139), .c(n138), .O(n141));
  or2    g0026(.a(n141), .b(n137), .O(n142));
  not    g0027(.a(in53), .O(n143));
  not    g0028(.a(in9), .O(n144));
  nand2  g0029(.a(n141), .b(n144), .O(n145));
  or2    g0030(.a(n145), .b(in78), .O(n146));
  not    g0031(.a(n146), .O(n147));
  nor3   g0032(.a(n147), .b(n143), .c(in49), .O(n148));
  xor2a  g0033(.a(n148), .b(n142), .O(n149));
  not    g0034(.a(n149), .O(n150));
  not    g0035(.a(in51), .O(n151));
  and2   g0036(.a(in98), .b(in24), .O(n152));
  not    g0037(.a(n152), .O(n153));
  xor2a  g0038(.a(in17), .b(in3), .O(n154));
  xor2a  g0039(.a(n154), .b(n127), .O(n155));
  and2   g0040(.a(n155), .b(n153), .O(n156));
  not    g0041(.a(n156), .O(n157));
  and2   g0042(.a(in106), .b(in23), .O(n158));
  or2    g0043(.a(n158), .b(n157), .O(n159));
  not    g0044(.a(n159), .O(n160));
  not    g0045(.a(in110), .O(n161));
  not    g0046(.a(in50), .O(n162));
  xor2a  g0047(.a(in64), .b(in40), .O(n163));
  xor2a  g0048(.a(n163), .b(in110), .O(n164));
  xnor2a g0049(.a(in84), .b(in52), .O(n165));
  xor2a  g0050(.a(n165), .b(n164), .O(n166));
  or2    g0051(.a(in110), .b(in73), .O(n167));
  not    g0052(.a(n142), .O(n168));
  nand4  g0053(.a(n168), .b(n167), .c(n166), .d(n162), .O(n169));
  nor2   g0054(.a(n169), .b(n155), .O(n170));
  not    g0055(.a(in63), .O(n171));
  not    g0056(.a(in30), .O(n172));
  xor2a  g0057(.a(in96), .b(in2), .O(n173));
  xor2a  g0058(.a(n173), .b(in51), .O(n174));
  xor2a  g0059(.a(n174), .b(n172), .O(n175));
  xor2a  g0060(.a(n175), .b(in112), .O(n176));
  xor2a  g0061(.a(in100), .b(in8), .O(n177));
  nor3   g0062(.a(n177), .b(in81), .c(in17), .O(n178));
  or2    g0063(.a(in85), .b(n131), .O(n179));
  or2    g0064(.a(n179), .b(n178), .O(n180));
  nand3  g0065(.a(n180), .b(n176), .c(n171), .O(n181));
  nand3  g0066(.a(n181), .b(n170), .c(n161), .O(n182));
  not    g0067(.a(n182), .O(n183));
  not    g0068(.a(in114), .O(n184));
  not    g0069(.a(in43), .O(n185));
  or2    g0070(.a(in60), .b(n185), .O(n186));
  xor2a  g0071(.a(n186), .b(n184), .O(n187));
  not    g0072(.a(in39), .O(n188));
  not    g0073(.a(in100), .O(n189));
  nand2  g0074(.a(n161), .b(n139), .O(n190));
  nand3  g0075(.a(n190), .b(n189), .c(n188), .O(n191));
  xor2a  g0076(.a(n191), .b(in90), .O(n192));
  not    g0077(.a(in16), .O(n193));
  nand3  g0078(.a(in104), .b(in48), .c(in28), .O(n194));
  nand3  g0079(.a(n194), .b(n141), .c(n138), .O(n195));
  xor2a  g0080(.a(n195), .b(n193), .O(n196));
  xor2a  g0081(.a(n196), .b(n192), .O(n197));
  not    g0082(.a(n197), .O(n198));
  not    g0083(.a(in69), .O(n199));
  not    g0084(.a(in56), .O(n200));
  not    g0085(.a(in68), .O(n201));
  not    g0086(.a(in70), .O(n202));
  nand4  g0087(.a(n202), .b(n201), .c(n200), .d(in50), .O(n203));
  xor2a  g0088(.a(n203), .b(n199), .O(n204));
  and2   g0089(.a(n204), .b(n155), .O(n205));
  nand3  g0090(.a(n205), .b(n198), .c(n187), .O(n206));
  not    g0091(.a(n206), .O(n207));
  nand4  g0092(.a(n207), .b(n183), .c(n160), .d(n151), .O(n208));
  xor2a  g0093(.a(n208), .b(n150), .O(n209));
  not    g0094(.a(n209), .O(n210));
  not    g0095(.a(in38), .O(n211));
  nor2   g0096(.a(n211), .b(in15), .O(n212));
  xor2a  g0097(.a(n145), .b(in91), .O(n213));
  xnor2a g0098(.a(n213), .b(n212), .O(n214));
  not    g0099(.a(in45), .O(n215));
  not    g0100(.a(in65), .O(n216));
  or2    g0101(.a(n216), .b(n215), .O(n217));
  and2   g0102(.a(in91), .b(in49), .O(n218));
  nand4  g0103(.a(in83), .b(in60), .c(in44), .d(in10), .O(n219));
  not    g0104(.a(n219), .O(n220));
  nand4  g0105(.a(n220), .b(n218), .c(n217), .d(in55), .O(n221));
  nand3  g0106(.a(n221), .b(n214), .c(n201), .O(n222));
  not    g0107(.a(n222), .O(n223));
  nand2  g0108(.a(n122), .b(n197), .O(n224));
  not    g0109(.a(in35), .O(n225));
  not    g0110(.a(in12), .O(n226));
  nand2  g0111(.a(in89), .b(in25), .O(n227));
  nand3  g0112(.a(n227), .b(n143), .c(n226), .O(n228));
  nand4  g0113(.a(n228), .b(in62), .c(in39), .d(n225), .O(n229));
  not    g0114(.a(n229), .O(n230));
  nand3  g0115(.a(n230), .b(n204), .c(n155), .O(n231));
  xor2a  g0116(.a(n231), .b(n215), .O(n232));
  xor2a  g0117(.a(n232), .b(n224), .O(n233));
  not    g0118(.a(in26), .O(n234));
  not    g0119(.a(in6), .O(n235));
  not    g0120(.a(in59), .O(n236));
  nand4  g0121(.a(in65), .b(n236), .c(in45), .d(n235), .O(n237));
  not    g0122(.a(in76), .O(n238));
  xor2a  g0123(.a(n227), .b(in30), .O(n239));
  nor2   g0124(.a(in98), .b(in18), .O(n240));
  nand3  g0125(.a(n240), .b(n239), .c(n238), .O(n241));
  not    g0126(.a(in32), .O(n242));
  xor2a  g0127(.a(in92), .b(in21), .O(n243));
  and2   g0128(.a(n243), .b(n242), .O(n244));
  xor2a  g0129(.a(in67), .b(in34), .O(n245));
  and2   g0130(.a(n245), .b(in9), .O(n246));
  nand4  g0131(.a(n246), .b(n244), .c(n241), .d(n237), .O(n247));
  nor3   g0132(.a(in113), .b(in74), .c(in17), .O(n248));
  or2    g0133(.a(in86), .b(in19), .O(n249));
  nor2   g0134(.a(n249), .b(n248), .O(n250));
  nand4  g0135(.a(n250), .b(in82), .c(in56), .d(n133), .O(n251));
  nor2   g0136(.a(n251), .b(n247), .O(n252));
  xor2a  g0137(.a(n252), .b(n234), .O(n253));
  nand2  g0138(.a(n253), .b(n233), .O(n254));
  xnor2a g0139(.a(n232), .b(n224), .O(n255));
  not    g0140(.a(n253), .O(n256));
  nand2  g0141(.a(n256), .b(n255), .O(n257));
  and2   g0142(.a(n159), .b(in114), .O(n258));
  nand3  g0143(.a(n258), .b(n257), .c(n254), .O(n259));
  nand2  g0144(.a(n259), .b(n223), .O(n260));
  nand3  g0145(.a(n192), .b(n177), .c(in50), .O(n261));
  not    g0146(.a(in108), .O(n262));
  and2   g0147(.a(n262), .b(in52), .O(n263));
  not    g0148(.a(in48), .O(n264));
  xor2a  g0149(.a(n142), .b(n264), .O(n265));
  xor2a  g0150(.a(n265), .b(n263), .O(n266));
  nand3  g0151(.a(n266), .b(n261), .c(in44), .O(n267));
  or2    g0152(.a(n267), .b(in35), .O(n268));
  not    g0153(.a(n268), .O(n269));
  nand2  g0154(.a(n269), .b(n260), .O(n270));
  nor3   g0155(.a(in111), .b(in66), .c(in17), .O(n271));
  xor2a  g0156(.a(n271), .b(in94), .O(n272));
  or2    g0157(.a(n272), .b(n204), .O(n273));
  xor2a  g0158(.a(n273), .b(in1), .O(n274));
  not    g0159(.a(n274), .O(n275));
  xor2a  g0160(.a(n275), .b(n270), .O(n276));
  not    g0161(.a(in27), .O(n277));
  not    g0162(.a(n187), .O(n278));
  not    g0163(.a(in77), .O(n279));
  or2    g0164(.a(n171), .b(in16), .O(n280));
  xor2a  g0165(.a(n280), .b(n279), .O(n281));
  xor2a  g0166(.a(n281), .b(n118), .O(n282));
  nand4  g0167(.a(n282), .b(n278), .c(in58), .d(n277), .O(n283));
  nand3  g0168(.a(in114), .b(in103), .c(in4), .O(n284));
  not    g0169(.a(n284), .O(n285));
  or2    g0170(.a(n285), .b(n143), .O(n286));
  nor2   g0171(.a(n286), .b(n283), .O(n287));
  and2   g0172(.a(in110), .b(in72), .O(n288));
  not    g0173(.a(n288), .O(n289));
  xor2a  g0174(.a(n289), .b(n287), .O(n290));
  xor2a  g0175(.a(n290), .b(n276), .O(n291));
  nand4  g0176(.a(n291), .b(n210), .c(n136), .d(n123), .O(n292));
  not    g0177(.a(in22), .O(n293));
  nand2  g0178(.a(in61), .b(n293), .O(n294));
  not    g0179(.a(in61), .O(n295));
  nand2  g0180(.a(n295), .b(in22), .O(n296));
  nand3  g0181(.a(n296), .b(n294), .c(in85), .O(n297));
  not    g0182(.a(in85), .O(n298));
  xor2a  g0183(.a(in61), .b(in22), .O(n299));
  nand2  g0184(.a(n299), .b(n298), .O(n300));
  nand3  g0185(.a(n300), .b(n297), .c(n215), .O(n301));
  not    g0186(.a(n301), .O(n302));
  nand3  g0187(.a(n300), .b(n297), .c(n162), .O(n303));
  xor2a  g0188(.a(n303), .b(in101), .O(n304));
  xor2a  g0189(.a(n304), .b(n302), .O(n305));
  nand2  g0190(.a(n305), .b(n180), .O(n306));
  not    g0191(.a(n180), .O(n307));
  xor2a  g0192(.a(n304), .b(n301), .O(n308));
  nand2  g0193(.a(n308), .b(n307), .O(n309));
  not    g0194(.a(in91), .O(n310));
  xnor2a g0195(.a(in99), .b(in13), .O(n311));
  xor2a  g0196(.a(in55), .b(in32), .O(n312));
  xor2a  g0197(.a(n312), .b(in36), .O(n313));
  not    g0198(.a(n313), .O(n314));
  nand3  g0199(.a(n314), .b(n311), .c(n310), .O(n315));
  not    g0200(.a(n315), .O(n316));
  nand3  g0201(.a(n316), .b(n309), .c(n306), .O(n317));
  xor2a  g0202(.a(n308), .b(n307), .O(n318));
  not    g0203(.a(n227), .O(n319));
  not    g0204(.a(in104), .O(n320));
  or2    g0205(.a(n219), .b(n320), .O(n321));
  or2    g0206(.a(n321), .b(n319), .O(n322));
  or2    g0207(.a(in88), .b(n151), .O(n323));
  xnor2a g0208(.a(n323), .b(in10), .O(n324));
  xor2a  g0209(.a(n324), .b(n322), .O(n325));
  nor2   g0210(.a(n325), .b(n157), .O(n326));
  nand4  g0211(.a(n326), .b(n316), .c(n318), .d(in107), .O(n327));
  and2   g0212(.a(n327), .b(n197), .O(n328));
  xor2a  g0213(.a(n328), .b(n317), .O(n329));
  xor2a  g0214(.a(n329), .b(in68), .O(n330));
  xor2a  g0215(.a(n330), .b(n292), .O(n331));
  not    g0216(.a(in29), .O(n332));
  not    g0217(.a(in99), .O(n333));
  nand4  g0218(.a(n262), .b(n333), .c(in52), .d(n332), .O(n334));
  not    g0219(.a(n334), .O(n335));
  not    g0220(.a(in37), .O(n336));
  xor2a  g0221(.a(n163), .b(n161), .O(n337));
  nand2  g0222(.a(n337), .b(n336), .O(n338));
  nand2  g0223(.a(n164), .b(in37), .O(n339));
  nand3  g0224(.a(n339), .b(n338), .c(n335), .O(n340));
  not    g0225(.a(n340), .O(n341));
  xor2a  g0226(.a(n213), .b(n212), .O(n342));
  xor2a  g0227(.a(n323), .b(n136), .O(n343));
  nand2  g0228(.a(n343), .b(n342), .O(n344));
  not    g0229(.a(in46), .O(n345));
  not    g0230(.a(in95), .O(n346));
  nand3  g0231(.a(n346), .b(n345), .c(in31), .O(n347));
  not    g0232(.a(n347), .O(n348));
  nand4  g0233(.a(in105), .b(in83), .c(in44), .d(in10), .O(n349));
  xor2a  g0234(.a(n349), .b(n235), .O(n350));
  xor2a  g0235(.a(n350), .b(n348), .O(n351));
  nand3  g0236(.a(n351), .b(n187), .c(n146), .O(n352));
  not    g0237(.a(n352), .O(n353));
  xor2a  g0238(.a(n353), .b(n344), .O(n354));
  or2    g0239(.a(n354), .b(n341), .O(n355));
  not    g0240(.a(in62), .O(n356));
  not    g0241(.a(n287), .O(n357));
  nand3  g0242(.a(n357), .b(n214), .c(n356), .O(n358));
  xor2a  g0243(.a(n358), .b(n355), .O(n359));
  not    g0244(.a(n359), .O(n360));
  xor2a  g0245(.a(n274), .b(n270), .O(n361));
  not    g0246(.a(in112), .O(n362));
  and2   g0247(.a(n273), .b(n160), .O(n363));
  not    g0248(.a(in84), .O(n364));
  xor2a  g0249(.a(in54), .b(in3), .O(n365));
  xor2a  g0250(.a(n365), .b(n364), .O(n366));
  not    g0251(.a(n366), .O(n367));
  not    g0252(.a(in78), .O(n368));
  nor2   g0253(.a(in110), .b(in58), .O(n369));
  nor2   g0254(.a(n369), .b(in109), .O(n370));
  xor2a  g0255(.a(n370), .b(n368), .O(n371));
  xor2a  g0256(.a(n371), .b(n129), .O(n372));
  xor2a  g0257(.a(n372), .b(n310), .O(n373));
  nand2  g0258(.a(n373), .b(n367), .O(n374));
  xor2a  g0259(.a(n372), .b(in91), .O(n375));
  nand2  g0260(.a(n375), .b(n366), .O(n376));
  nand4  g0261(.a(n376), .b(n374), .c(n284), .d(in40), .O(n377));
  nand3  g0262(.a(n377), .b(n122), .c(n223), .O(n378));
  and2   g0263(.a(n342), .b(in93), .O(n379));
  nand3  g0264(.a(n379), .b(n378), .c(n221), .O(n380));
  xor2a  g0265(.a(n380), .b(n363), .O(n381));
  not    g0266(.a(n381), .O(n382));
  xor2a  g0267(.a(n212), .b(n171), .O(n383));
  xor2a  g0268(.a(n383), .b(n222), .O(n384));
  xor2a  g0269(.a(n384), .b(n317), .O(n385));
  xor2a  g0270(.a(n381), .b(n385), .O(n386));
  not    g0271(.a(n252), .O(n387));
  and2   g0272(.a(n387), .b(in20), .O(n388));
  xor2a  g0273(.a(n288), .b(n247), .O(n389));
  not    g0274(.a(n311), .O(n390));
  or2    g0275(.a(n313), .b(n390), .O(n391));
  nand2  g0276(.a(n283), .b(n391), .O(n392));
  xnor2a g0277(.a(in79), .b(in78), .O(n393));
  xnor2a g0278(.a(n393), .b(n392), .O(n394));
  nand3  g0279(.a(n394), .b(n389), .c(n116), .O(n395));
  and2   g0280(.a(n395), .b(n347), .O(n396));
  nor2   g0281(.a(n396), .b(in9), .O(n397));
  and2   g0282(.a(n270), .b(n236), .O(n398));
  nand4  g0283(.a(n398), .b(n397), .c(n388), .d(n386), .O(n399));
  nand2  g0284(.a(n399), .b(n354), .O(n400));
  or2    g0285(.a(in111), .b(in57), .O(n401));
  xnor2a g0286(.a(n271), .b(n135), .O(n402));
  nand3  g0287(.a(n314), .b(n311), .c(n263), .O(n403));
  xnor2a g0288(.a(n403), .b(n402), .O(n404));
  xor2a  g0289(.a(n285), .b(n243), .O(n405));
  xnor2a g0290(.a(n405), .b(n404), .O(n406));
  not    g0291(.a(n406), .O(n407));
  nor4   g0292(.a(n267), .b(n407), .c(n221), .d(n184), .O(n408));
  xor2a  g0293(.a(n408), .b(n401), .O(n409));
  xor2a  g0294(.a(n409), .b(n400), .O(n410));
  nand2  g0295(.a(n410), .b(n382), .O(n411));
  not    g0296(.a(in47), .O(n412));
  not    g0297(.a(n135), .O(n413));
  not    g0298(.a(in81), .O(n414));
  and2   g0299(.a(in95), .b(n414), .O(n415));
  nand4  g0300(.a(n415), .b(n314), .c(n413), .d(n226), .O(n416));
  not    g0301(.a(n416), .O(n417));
  nor3   g0302(.a(n417), .b(in69), .c(n412), .O(n418));
  nand3  g0303(.a(n244), .b(n241), .c(n237), .O(n419));
  not    g0304(.a(n349), .O(n420));
  nand4  g0305(.a(n220), .b(n420), .c(in104), .d(n414), .O(n421));
  not    g0306(.a(n421), .O(n422));
  nand4  g0307(.a(n422), .b(n402), .c(n419), .d(n117), .O(n423));
  not    g0308(.a(in28), .O(n424));
  not    g0309(.a(n165), .O(n425));
  nand3  g0310(.a(n401), .b(n425), .c(n424), .O(n426));
  xor2a  g0311(.a(n288), .b(n426), .O(n427));
  xor2a  g0312(.a(n427), .b(n423), .O(n428));
  xor2a  g0313(.a(n428), .b(in111), .O(n429));
  xor2a  g0314(.a(n429), .b(n287), .O(n430));
  nor3   g0315(.a(n313), .b(in107), .c(in53), .O(n431));
  or2    g0316(.a(n431), .b(n168), .O(n432));
  not    g0317(.a(in82), .O(n433));
  and2   g0318(.a(n152), .b(n433), .O(n434));
  nand3  g0319(.a(n421), .b(n289), .c(in9), .O(n435));
  nand4  g0320(.a(n435), .b(n434), .c(n432), .d(in99), .O(n436));
  not    g0321(.a(n436), .O(n437));
  nand4  g0322(.a(n437), .b(n430), .c(n418), .d(in107), .O(n438));
  nand2  g0323(.a(n209), .b(n279), .O(n439));
  nor2   g0324(.a(n439), .b(n438), .O(n440));
  not    g0325(.a(n440), .O(n441));
  nand3  g0326(.a(n402), .b(n419), .c(n117), .O(n442));
  not    g0327(.a(n442), .O(n443));
  and2   g0328(.a(n244), .b(n241), .O(n444));
  not    g0329(.a(in20), .O(n445));
  nand3  g0330(.a(n342), .b(n341), .c(in38), .O(n446));
  xor2a  g0331(.a(n446), .b(n445), .O(n447));
  nand4  g0332(.a(n447), .b(n156), .c(n444), .d(in94), .O(n448));
  nand3  g0333(.a(n156), .b(n444), .c(in94), .O(n449));
  xor2a  g0334(.a(n446), .b(in20), .O(n450));
  nand2  g0335(.a(n450), .b(n449), .O(n451));
  not    g0336(.a(in89), .O(n452));
  nand3  g0337(.a(n403), .b(n452), .c(in69), .O(n453));
  or2    g0338(.a(n453), .b(n295), .O(n454));
  not    g0339(.a(n454), .O(n455));
  xor2a  g0340(.a(n152), .b(n445), .O(n456));
  not    g0341(.a(n228), .O(n457));
  nor3   g0342(.a(n457), .b(n356), .c(n188), .O(n458));
  nand4  g0343(.a(n458), .b(n456), .c(n166), .d(n277), .O(n459));
  not    g0344(.a(n459), .O(n460));
  and2   g0345(.a(n460), .b(n211), .O(n461));
  nand4  g0346(.a(n461), .b(n455), .c(n451), .d(n448), .O(n462));
  nand2  g0347(.a(n462), .b(n443), .O(n463));
  xor2a  g0348(.a(n463), .b(n278), .O(n464));
  xor2a  g0349(.a(in108), .b(in51), .O(n465));
  xor2a  g0350(.a(n303), .b(in26), .O(n466));
  xor2a  g0351(.a(n466), .b(n465), .O(n467));
  not    g0352(.a(n322), .O(n468));
  nand4  g0353(.a(n468), .b(n316), .c(n318), .d(in71), .O(n469));
  nand2  g0354(.a(n469), .b(n160), .O(n470));
  and2   g0355(.a(n470), .b(n467), .O(n471));
  xor2a  g0356(.a(n259), .b(in55), .O(n472));
  xor2a  g0357(.a(n472), .b(n471), .O(n473));
  xor2a  g0358(.a(n473), .b(n424), .O(n474));
  nand2  g0359(.a(n474), .b(n464), .O(n475));
  not    g0360(.a(n464), .O(n476));
  xor2a  g0361(.a(n473), .b(in28), .O(n477));
  nand2  g0362(.a(n477), .b(n476), .O(n478));
  nand4  g0363(.a(n478), .b(n475), .c(n441), .d(n352), .O(n479));
  not    g0364(.a(n479), .O(n480));
  nand3  g0365(.a(n480), .b(n411), .c(n362), .O(n481));
  nand2  g0366(.a(n481), .b(n361), .O(n482));
  or2    g0367(.a(n359), .b(n366), .O(n483));
  not    g0368(.a(n328), .O(n484));
  not    g0369(.a(n205), .O(n485));
  nand3  g0370(.a(n273), .b(n485), .c(n264), .O(n486));
  xor2a  g0371(.a(n204), .b(in89), .O(n487));
  xor2a  g0372(.a(n487), .b(n486), .O(n488));
  and2   g0373(.a(n488), .b(n363), .O(n489));
  xor2a  g0374(.a(n385), .b(n404), .O(n490));
  nand3  g0375(.a(n301), .b(n320), .c(n234), .O(n491));
  xor2a  g0376(.a(n135), .b(in71), .O(n492));
  xor2a  g0377(.a(n492), .b(n491), .O(n493));
  nand3  g0378(.a(n493), .b(n186), .c(in39), .O(n494));
  not    g0379(.a(n494), .O(n495));
  not    g0380(.a(in33), .O(n496));
  nand2  g0381(.a(n240), .b(n239), .O(n497));
  not    g0382(.a(n497), .O(n498));
  and2   g0383(.a(n202), .b(in11), .O(n499));
  or2    g0384(.a(n499), .b(in47), .O(n500));
  nand3  g0385(.a(n500), .b(n498), .c(n215), .O(n501));
  xor2a  g0386(.a(n501), .b(in18), .O(n502));
  xor2a  g0387(.a(n502), .b(n496), .O(n503));
  xor2a  g0388(.a(n503), .b(n436), .O(n504));
  xor2a  g0389(.a(n504), .b(n421), .O(n505));
  xor2a  g0390(.a(n214), .b(in8), .O(n506));
  xor2a  g0391(.a(n506), .b(n505), .O(n507));
  nand2  g0392(.a(n507), .b(n495), .O(n508));
  nand3  g0393(.a(n473), .b(n508), .c(in90), .O(n509));
  nand3  g0394(.a(n509), .b(n490), .c(in38), .O(n510));
  not    g0395(.a(n510), .O(n511));
  nand3  g0396(.a(n511), .b(n489), .c(in56), .O(n512));
  not    g0397(.a(n247), .O(n513));
  nand3  g0398(.a(n181), .b(n513), .c(n141), .O(n514));
  not    g0399(.a(n514), .O(n515));
  nand4  g0400(.a(n360), .b(n515), .c(n367), .d(n264), .O(n516));
  nand4  g0401(.a(n516), .b(n378), .c(n489), .d(in59), .O(n517));
  xnor2a g0402(.a(n517), .b(n510), .O(n518));
  nand3  g0403(.a(n518), .b(n512), .c(n117), .O(n519));
  or2    g0404(.a(n519), .b(n484), .O(n520));
  or2    g0405(.a(n520), .b(n483), .O(n521));
  and2   g0406(.a(n521), .b(n252), .O(n522));
  not    g0407(.a(n191), .O(n523));
  and2   g0408(.a(in83), .b(in10), .O(n524));
  not    g0409(.a(in102), .O(n525));
  and2   g0410(.a(n497), .b(n525), .O(n526));
  xnor2a g0411(.a(n526), .b(n141), .O(n527));
  xnor2a g0412(.a(n467), .b(n241), .O(n528));
  xnor2a g0413(.a(in87), .b(in61), .O(n529));
  xor2a  g0414(.a(n529), .b(n177), .O(n530));
  xor2a  g0415(.a(n530), .b(n528), .O(n531));
  and2   g0416(.a(n342), .b(in114), .O(n532));
  nand4  g0417(.a(n532), .b(n531), .c(n148), .d(n527), .O(n533));
  not    g0418(.a(in72), .O(n534));
  and2   g0419(.a(n389), .b(n534), .O(n535));
  nand4  g0420(.a(n535), .b(n357), .c(n326), .d(n390), .O(n536));
  and2   g0421(.a(n536), .b(n495), .O(n537));
  xor2a  g0422(.a(n537), .b(n533), .O(n538));
  not    g0423(.a(n438), .O(n539));
  nor3   g0424(.a(n539), .b(n538), .c(n120), .O(n540));
  nor3   g0425(.a(n206), .b(n540), .c(n524), .O(n541));
  nand2  g0426(.a(n377), .b(n193), .O(n542));
  nor2   g0427(.a(n542), .b(n209), .O(n543));
  not    g0428(.a(in66), .O(n544));
  and2   g0429(.a(n247), .b(in13), .O(n545));
  not    g0430(.a(n145), .O(n546));
  not    g0431(.a(in3), .O(n547));
  xnor2a g0432(.a(in103), .b(in19), .O(n548));
  or2    g0433(.a(n548), .b(n184), .O(n549));
  xor2a  g0434(.a(n549), .b(n547), .O(n550));
  xor2a  g0435(.a(n550), .b(n546), .O(n551));
  xor2a  g0436(.a(n191), .b(in72), .O(n552));
  xor2a  g0437(.a(n552), .b(n178), .O(n553));
  nand3  g0438(.a(n553), .b(n551), .c(in85), .O(n554));
  nand4  g0439(.a(n554), .b(n178), .c(n545), .d(n527), .O(n555));
  not    g0440(.a(in79), .O(n556));
  not    g0441(.a(in4), .O(n557));
  xor2a  g0442(.a(n494), .b(n557), .O(n558));
  xor2a  g0443(.a(n558), .b(n406), .O(n559));
  nand2  g0444(.a(n559), .b(n556), .O(n560));
  nand2  g0445(.a(n560), .b(n153), .O(n561));
  nand3  g0446(.a(n561), .b(n555), .c(n544), .O(n562));
  xor2a  g0447(.a(n562), .b(n543), .O(n563));
  nand2  g0448(.a(n563), .b(n508), .O(n564));
  nand3  g0449(.a(n564), .b(n252), .c(in30), .O(n565));
  nor4   g0450(.a(n565), .b(n541), .c(n170), .d(n414), .O(n566));
  not    g0451(.a(in94), .O(n567));
  nand2  g0452(.a(n528), .b(in80), .O(n568));
  xor2a  g0453(.a(n528), .b(in87), .O(n569));
  xor2a  g0454(.a(n569), .b(n568), .O(n570));
  not    g0455(.a(in25), .O(n571));
  xor2a  g0456(.a(n432), .b(n242), .O(n572));
  xor2a  g0457(.a(n572), .b(n252), .O(n573));
  nand3  g0458(.a(n462), .b(n573), .c(n571), .O(n574));
  nand3  g0459(.a(n574), .b(n570), .c(n567), .O(n575));
  or2    g0460(.a(n394), .b(n424), .O(n576));
  not    g0461(.a(n576), .O(n577));
  nand4  g0462(.a(n577), .b(n464), .c(n575), .d(in84), .O(n578));
  nand2  g0463(.a(n290), .b(n276), .O(n579));
  not    g0464(.a(n290), .O(n580));
  nand2  g0465(.a(n580), .b(n361), .O(n581));
  nand4  g0466(.a(n581), .b(n579), .c(n578), .d(in10), .O(n582));
  nand3  g0467(.a(n582), .b(n564), .c(in65), .O(n583));
  nand2  g0468(.a(n583), .b(n385), .O(n584));
  and2   g0469(.a(n555), .b(n459), .O(n585));
  xor2a  g0470(.a(n585), .b(n355), .O(n586));
  nor2   g0471(.a(n586), .b(n557), .O(n587));
  nand2  g0472(.a(n587), .b(n584), .O(n588));
  xor2a  g0473(.a(n471), .b(n225), .O(n589));
  xor2a  g0474(.a(n589), .b(n588), .O(n590));
  nand3  g0475(.a(n590), .b(n566), .c(in63), .O(n591));
  nand3  g0476(.a(n509), .b(n591), .c(n523), .O(n592));
  xor2a  g0477(.a(n592), .b(in101), .O(n593));
  xor2a  g0478(.a(n593), .b(n522), .O(n594));
  not    g0479(.a(n594), .O(n595));
  or2    g0480(.a(n595), .b(n387), .O(n596));
  nand3  g0481(.a(n397), .b(n388), .c(n386), .O(n597));
  not    g0482(.a(n597), .O(n598));
  not    g0483(.a(n354), .O(n599));
  or2    g0484(.a(n197), .b(n278), .O(n600));
  nand4  g0485(.a(n395), .b(n600), .c(n347), .d(in81), .O(n601));
  xor2a  g0486(.a(n601), .b(n209), .O(n602));
  xor2a  g0487(.a(n602), .b(n159), .O(n603));
  or2    g0488(.a(n603), .b(n599), .O(n604));
  nand2  g0489(.a(n604), .b(n267), .O(n605));
  xor2a  g0490(.a(n509), .b(n547), .O(n606));
  xor2a  g0491(.a(n606), .b(n605), .O(n607));
  nand3  g0492(.a(n607), .b(n331), .c(n361), .O(n608));
  not    g0493(.a(n329), .O(n609));
  xnor2a g0494(.a(n149), .b(in52), .O(n610));
  xor2a  g0495(.a(n610), .b(n440), .O(n611));
  xor2a  g0496(.a(n570), .b(in81), .O(n612));
  xor2a  g0497(.a(n612), .b(n611), .O(n613));
  nand3  g0498(.a(n613), .b(n259), .c(n119), .O(n614));
  nand3  g0499(.a(n614), .b(n609), .c(in113), .O(n615));
  not    g0500(.a(n291), .O(n616));
  and2   g0501(.a(n616), .b(n445), .O(n617));
  not    g0502(.a(n273), .O(n618));
  or2    g0503(.a(n618), .b(in3), .O(n619));
  nor4   g0504(.a(n619), .b(n267), .c(n149), .d(n144), .O(n620));
  xor2a  g0505(.a(n260), .b(n140), .O(n621));
  xor2a  g0506(.a(n621), .b(n620), .O(n622));
  nand3  g0507(.a(n622), .b(n210), .c(n271), .O(n623));
  nand2  g0508(.a(n623), .b(n509), .O(n624));
  xor2a  g0509(.a(n327), .b(in43), .O(n625));
  xor2a  g0510(.a(n625), .b(n624), .O(n626));
  xor2a  g0511(.a(n626), .b(n469), .O(n627));
  nand4  g0512(.a(n627), .b(n617), .c(n615), .d(n370), .O(n628));
  not    g0513(.a(n395), .O(n629));
  nand4  g0514(.a(n511), .b(n380), .c(n489), .d(in56), .O(n630));
  nand2  g0515(.a(n630), .b(n480), .O(n631));
  not    g0516(.a(n426), .O(n632));
  or2    g0517(.a(n632), .b(n459), .O(n633));
  xor2a  g0518(.a(n633), .b(n570), .O(n634));
  or2    g0519(.a(n182), .b(n390), .O(n635));
  not    g0520(.a(n635), .O(n636));
  and2   g0521(.a(n636), .b(n634), .O(n637));
  xor2a  g0522(.a(n637), .b(in57), .O(n638));
  xor2a  g0523(.a(n638), .b(n631), .O(n639));
  not    g0524(.a(n503), .O(n640));
  nor2   g0525(.a(n640), .b(n533), .O(n641));
  xor2a  g0526(.a(n490), .b(n364), .O(n642));
  xor2a  g0527(.a(n642), .b(n641), .O(n643));
  xor2a  g0528(.a(n643), .b(n129), .O(n644));
  xor2a  g0529(.a(n644), .b(n639), .O(n645));
  nand3  g0530(.a(n645), .b(n629), .c(n473), .O(n646));
  and2   g0531(.a(n533), .b(n413), .O(n647));
  or2    g0532(.a(n616), .b(in70), .O(n648));
  not    g0533(.a(n648), .O(n649));
  nand4  g0534(.a(n649), .b(n647), .c(n646), .d(n598), .O(n650));
  or2    g0535(.a(n536), .b(n158), .O(n651));
  nor2   g0536(.a(n651), .b(n650), .O(n652));
  nand2  g0537(.a(n388), .b(n386), .O(n653));
  xor2a  g0538(.a(n653), .b(n412), .O(n654));
  xor2a  g0539(.a(n654), .b(n652), .O(n655));
  nand2  g0540(.a(n655), .b(n628), .O(n656));
  nand3  g0541(.a(n656), .b(n464), .c(in113), .O(n657));
  not    g0542(.a(n260), .O(n658));
  not    g0543(.a(in107), .O(n659));
  nand4  g0544(.a(n636), .b(n634), .c(n354), .d(n525), .O(n660));
  or2    g0545(.a(n660), .b(n460), .O(n661));
  not    g0546(.a(n661), .O(n662));
  nand3  g0547(.a(n662), .b(n660), .c(n659), .O(n663));
  and2   g0548(.a(n663), .b(n658), .O(n664));
  or2    g0549(.a(n430), .b(n664), .O(n665));
  not    g0550(.a(in36), .O(n666));
  xor2a  g0551(.a(n359), .b(n666), .O(n667));
  xor2a  g0552(.a(n667), .b(n665), .O(n668));
  xor2a  g0553(.a(n668), .b(n361), .O(n669));
  xor2a  g0554(.a(n669), .b(n179), .O(n670));
  xor2a  g0555(.a(n670), .b(n657), .O(n671));
  nand2  g0556(.a(n671), .b(n608), .O(n672));
  and2   g0557(.a(n653), .b(n184), .O(n673));
  and2   g0558(.a(n614), .b(n321), .O(n674));
  nand3  g0559(.a(n674), .b(n673), .c(n672), .O(n675));
  not    g0560(.a(n453), .O(n676));
  not    g0561(.a(n380), .O(n677));
  nand2  g0562(.a(n586), .b(n546), .O(n678));
  xor2a  g0563(.a(n447), .b(n449), .O(n679));
  xor2a  g0564(.a(n679), .b(in19), .O(n680));
  xnor2a g0565(.a(n680), .b(n678), .O(n681));
  nand3  g0566(.a(n681), .b(n677), .c(in98), .O(n682));
  nand3  g0567(.a(n250), .b(in82), .c(in56), .O(n683));
  not    g0568(.a(n683), .O(n684));
  or2    g0569(.a(n514), .b(n149), .O(n685));
  nand3  g0570(.a(n685), .b(n392), .c(n684), .O(n686));
  or2    g0571(.a(n260), .b(n364), .O(n687));
  not    g0572(.a(n687), .O(n688));
  nand2  g0573(.a(n688), .b(n643), .O(n689));
  nand2  g0574(.a(n689), .b(n686), .O(n690));
  xor2a  g0575(.a(n690), .b(n666), .O(n691));
  xor2a  g0576(.a(n691), .b(n682), .O(n692));
  nand3  g0577(.a(n478), .b(n475), .c(n441), .O(n693));
  or2    g0578(.a(n693), .b(n567), .O(n694));
  not    g0579(.a(n694), .O(n695));
  nand2  g0580(.a(n695), .b(n692), .O(n696));
  nand3  g0581(.a(n617), .b(n615), .c(in62), .O(n697));
  not    g0582(.a(n697), .O(n698));
  nand3  g0583(.a(n698), .b(n696), .c(n608), .O(n699));
  nand2  g0584(.a(n699), .b(n676), .O(n700));
  not    g0585(.a(n512), .O(n701));
  nand2  g0586(.a(n589), .b(n588), .O(n702));
  not    g0587(.a(n589), .O(n703));
  nand3  g0588(.a(n703), .b(n587), .c(n584), .O(n704));
  nand3  g0589(.a(n704), .b(n702), .c(n209), .O(n705));
  xor2a  g0590(.a(n705), .b(n486), .O(n706));
  nand2  g0591(.a(n706), .b(n701), .O(n707));
  not    g0592(.a(n486), .O(n708));
  xor2a  g0593(.a(n705), .b(n708), .O(n709));
  nand2  g0594(.a(n709), .b(n512), .O(n710));
  nand4  g0595(.a(n710), .b(n707), .c(n700), .d(n234), .O(n711));
  not    g0596(.a(in17), .O(n712));
  and2   g0597(.a(n693), .b(n712), .O(n713));
  nand2  g0598(.a(n713), .b(n711), .O(n714));
  nand2  g0599(.a(n714), .b(n633), .O(n715));
  xor2a  g0600(.a(n715), .b(n663), .O(n716));
  xor2a  g0601(.a(n716), .b(in108), .O(n717));
  xnor2a g0602(.a(n717), .b(n675), .O(n718));
  or2    g0603(.a(n718), .b(n562), .O(n719));
  xor2a  g0604(.a(n719), .b(n598), .O(n720));
  or2    g0605(.a(n720), .b(n596), .O(n721));
  not    g0606(.a(n721), .O(n722));
  or2    g0607(.a(n722), .b(n479), .O(n723));
  nand2  g0608(.a(n723), .b(n482), .O(n724));
  xor2a  g0609(.a(n724), .b(n360), .O(n725));
  not    g0610(.a(n614), .O(n726));
  not    g0611(.a(n326), .O(n727));
  not    g0612(.a(n408), .O(n728));
  nand2  g0613(.a(n545), .b(n527), .O(n729));
  and2   g0614(.a(n729), .b(in103), .O(n730));
  nand4  g0615(.a(n730), .b(n728), .c(n209), .d(in57), .O(n731));
  xor2a  g0616(.a(n469), .b(n137), .O(n732));
  xor2a  g0617(.a(n732), .b(n731), .O(n733));
  nand2  g0618(.a(n733), .b(n153), .O(n734));
  nor2   g0619(.a(n734), .b(n512), .O(n735));
  not    g0620(.a(n490), .O(n736));
  or2    g0621(.a(n416), .b(n736), .O(n737));
  nand3  g0622(.a(n484), .b(n737), .c(n401), .O(n738));
  xnor2a g0623(.a(n738), .b(n686), .O(n739));
  xor2a  g0624(.a(n259), .b(n666), .O(n740));
  xnor2a g0625(.a(n740), .b(n739), .O(n741));
  nand2  g0626(.a(n741), .b(n735), .O(n742));
  nand2  g0627(.a(n742), .b(n727), .O(n743));
  xor2a  g0628(.a(n543), .b(n666), .O(n744));
  xor2a  g0629(.a(n744), .b(n743), .O(n745));
  nand2  g0630(.a(n745), .b(n538), .O(n746));
  not    g0631(.a(n746), .O(n747));
  and2   g0632(.a(n516), .b(in97), .O(n748));
  nand4  g0633(.a(n748), .b(n681), .c(n747), .d(in92), .O(n749));
  nand4  g0634(.a(n749), .b(n726), .c(n436), .d(n336), .O(n750));
  nand3  g0635(.a(n750), .b(n725), .c(n199), .O(n751));
  nand2  g0636(.a(n608), .b(n735), .O(n752));
  nand3  g0637(.a(n752), .b(n462), .c(n132), .O(n753));
  xnor2a g0638(.a(n753), .b(in40), .O(n754));
  xor2a  g0639(.a(n754), .b(n751), .O(n755));
  or2    g0640(.a(n755), .b(n331), .O(n756));
  not    g0641(.a(n756), .O(n757));
  nand3  g0642(.a(n663), .b(n658), .c(in18), .O(n758));
  not    g0643(.a(n758), .O(n759));
  and2   g0644(.a(n759), .b(n592), .O(n760));
  not    g0645(.a(in74), .O(n761));
  and2   g0646(.a(n736), .b(n761), .O(n762));
  nand3  g0647(.a(n762), .b(n481), .c(n361), .O(n763));
  not    g0648(.a(in57), .O(n764));
  and2   g0649(.a(n598), .b(n764), .O(n765));
  nand2  g0650(.a(n765), .b(n763), .O(n766));
  xor2a  g0651(.a(n366), .b(n678), .O(n767));
  not    g0652(.a(n767), .O(n768));
  xor2a  g0653(.a(n768), .b(n766), .O(n769));
  xor2a  g0654(.a(n400), .b(in46), .O(n770));
  xor2a  g0655(.a(n770), .b(n769), .O(n771));
  nand2  g0656(.a(n771), .b(n760), .O(n772));
  nand2  g0657(.a(n772), .b(n489), .O(n773));
  xor2a  g0658(.a(n746), .b(n263), .O(n774));
  xor2a  g0659(.a(n774), .b(n773), .O(n775));
  xor2a  g0660(.a(n741), .b(in17), .O(n776));
  xor2a  g0661(.a(n776), .b(n775), .O(n777));
  not    g0662(.a(n578), .O(n778));
  and2   g0663(.a(n778), .b(in36), .O(n779));
  or2    g0664(.a(n773), .b(n137), .O(n780));
  not    g0665(.a(n780), .O(n781));
  nand3  g0666(.a(n781), .b(n779), .c(n777), .O(n782));
  and2   g0667(.a(n563), .b(in77), .O(n783));
  and2   g0668(.a(n783), .b(n782), .O(n784));
  nand3  g0669(.a(n430), .b(n418), .c(in107), .O(n785));
  not    g0670(.a(n483), .O(n786));
  not    g0671(.a(n663), .O(n787));
  nand3  g0672(.a(n714), .b(n787), .c(n633), .O(n788));
  nand2  g0673(.a(n715), .b(n663), .O(n789));
  and2   g0674(.a(n689), .b(n158), .O(n790));
  nand3  g0675(.a(n790), .b(n789), .c(n788), .O(n791));
  nand2  g0676(.a(n791), .b(n585), .O(n792));
  not    g0677(.a(n585), .O(n793));
  nand4  g0678(.a(n790), .b(n789), .c(n788), .d(n793), .O(n794));
  and2   g0679(.a(n653), .b(n632), .O(n795));
  nand3  g0680(.a(n795), .b(n794), .c(n792), .O(n796));
  xor2a  g0681(.a(n737), .b(n304), .O(n797));
  xor2a  g0682(.a(n797), .b(n796), .O(n798));
  xor2a  g0683(.a(n798), .b(n786), .O(n799));
  nand2  g0684(.a(n799), .b(n785), .O(n800));
  xor2a  g0685(.a(n749), .b(n523), .O(n801));
  xor2a  g0686(.a(n801), .b(n800), .O(n802));
  nand2  g0687(.a(n802), .b(n733), .O(n803));
  not    g0688(.a(n208), .O(n804));
  not    g0689(.a(n627), .O(n805));
  nand4  g0690(.a(n613), .b(n480), .c(n140), .d(n764), .O(n806));
  nand4  g0691(.a(n806), .b(n515), .c(n150), .d(in9), .O(n807));
  nand3  g0692(.a(n807), .b(n805), .c(n727), .O(n808));
  nand3  g0693(.a(n783), .b(n782), .c(n207), .O(n809));
  nand2  g0694(.a(n809), .b(n808), .O(n810));
  and2   g0695(.a(n773), .b(n137), .O(n811));
  nand2  g0696(.a(n811), .b(n810), .O(n812));
  xor2a  g0697(.a(n812), .b(n489), .O(n813));
  xor2a  g0698(.a(n813), .b(n804), .O(n814));
  xor2a  g0699(.a(n623), .b(in83), .O(n815));
  xor2a  g0700(.a(n815), .b(n814), .O(n816));
  nand2  g0701(.a(n218), .b(n217), .O(n817));
  xor2a  g0702(.a(n540), .b(n817), .O(n818));
  not    g0703(.a(n818), .O(n819));
  xor2a  g0704(.a(n819), .b(n816), .O(n820));
  nand3  g0705(.a(n647), .b(n646), .c(n598), .O(n821));
  xor2a  g0706(.a(n821), .b(n203), .O(n822));
  nand2  g0707(.a(n822), .b(n820), .O(n823));
  xor2a  g0708(.a(n818), .b(n816), .O(n824));
  not    g0709(.a(n822), .O(n825));
  nand2  g0710(.a(n825), .b(n824), .O(n826));
  or2    g0711(.a(n520), .b(in31), .O(n827));
  not    g0712(.a(n827), .O(n828));
  nand3  g0713(.a(n828), .b(n826), .c(n823), .O(n829));
  xor2a  g0714(.a(n829), .b(n803), .O(n830));
  xor2a  g0715(.a(n830), .b(n471), .O(n831));
  xor2a  g0716(.a(n831), .b(n784), .O(n832));
  xor2a  g0717(.a(n363), .b(n194), .O(n833));
  xor2a  g0718(.a(n833), .b(n628), .O(n834));
  xor2a  g0719(.a(n743), .b(in47), .O(n835));
  xor2a  g0720(.a(n835), .b(n834), .O(n836));
  nand3  g0721(.a(n836), .b(n692), .c(in93), .O(n837));
  xor2a  g0722(.a(n837), .b(n753), .O(n838));
  xor2a  g0723(.a(n641), .b(n302), .O(n839));
  xor2a  g0724(.a(n839), .b(n838), .O(n840));
  xor2a  g0725(.a(n570), .b(n556), .O(n841));
  xor2a  g0726(.a(n841), .b(n808), .O(n842));
  xor2a  g0727(.a(n842), .b(in97), .O(n843));
  xor2a  g0728(.a(n843), .b(n840), .O(n844));
  not    g0729(.a(n844), .O(n845));
  or2    g0730(.a(n845), .b(n368), .O(n846));
  not    g0731(.a(n846), .O(n847));
  nand2  g0732(.a(n847), .b(n832), .O(n848));
  xor2a  g0733(.a(n650), .b(n320), .O(n849));
  xor2a  g0734(.a(n849), .b(n848), .O(n850));
  nand2  g0735(.a(n850), .b(n490), .O(n851));
  not    g0736(.a(n536), .O(n852));
  nand2  g0737(.a(n673), .b(n672), .O(n853));
  xor2a  g0738(.a(n657), .b(n735), .O(n854));
  xor2a  g0739(.a(n854), .b(n678), .O(n855));
  and2   g0740(.a(n855), .b(n853), .O(n856));
  nand3  g0741(.a(n718), .b(n856), .c(n199), .O(n857));
  xor2a  g0742(.a(n749), .b(in98), .O(n858));
  xor2a  g0743(.a(n858), .b(n857), .O(n859));
  xor2a  g0744(.a(n859), .b(n852), .O(n860));
  xor2a  g0745(.a(n860), .b(n681), .O(n861));
  xor2a  g0746(.a(n861), .b(in37), .O(n862));
  xor2a  g0747(.a(n862), .b(n851), .O(n863));
  nand2  g0748(.a(n863), .b(n664), .O(n864));
  nor2   g0749(.a(n856), .b(n456), .O(n865));
  nand2  g0750(.a(n865), .b(n864), .O(n866));
  not    g0751(.a(n462), .O(n867));
  xor2a  g0752(.a(n803), .b(n867), .O(n868));
  xor2a  g0753(.a(n868), .b(n785), .O(n869));
  or2    g0754(.a(n745), .b(in13), .O(n870));
  not    g0755(.a(n870), .O(n871));
  nand2  g0756(.a(n871), .b(n869), .O(n872));
  xor2a  g0757(.a(n756), .b(n653), .O(n873));
  nand2  g0758(.a(n872), .b(n844), .O(n874));
  nand2  g0759(.a(n874), .b(n793), .O(n875));
  xnor2a g0760(.a(n875), .b(n167), .O(n876));
  xor2a  g0761(.a(n876), .b(n873), .O(n877));
  nand2  g0762(.a(n877), .b(n872), .O(n878));
  nand2  g0763(.a(n878), .b(n866), .O(n879));
  nor2   g0764(.a(n631), .b(n348), .O(n880));
  nand4  g0765(.a(n880), .b(n879), .c(n586), .d(n546), .O(n881));
  xnor2a g0766(.a(n753), .b(n266), .O(n882));
  xor2a  g0767(.a(n882), .b(n881), .O(n883));
  xor2a  g0768(.a(n856), .b(in91), .O(n884));
  xor2a  g0769(.a(n884), .b(n883), .O(n885));
  nand3  g0770(.a(n885), .b(n757), .c(n122), .O(n886));
  xor2a  g0771(.a(n522), .b(in84), .O(n887));
  not    g0772(.a(n887), .O(n888));
  xor2a  g0773(.a(n888), .b(n886), .O(n889));
  not    g0774(.a(n889), .O(n890));
  not    g0775(.a(n583), .O(n891));
  not    g0776(.a(n874), .O(n892));
  nand2  g0777(.a(n892), .b(n866), .O(n893));
  nand2  g0778(.a(n893), .b(n745), .O(n894));
  nand2  g0779(.a(n894), .b(n891), .O(n895));
  nand3  g0780(.a(n893), .b(n745), .c(n583), .O(n896));
  not    g0781(.a(n615), .O(n897));
  not    g0782(.a(n126), .O(n898));
  not    g0783(.a(n696), .O(n899));
  nand4  g0784(.a(n594), .b(n899), .c(n252), .d(n898), .O(n900));
  nand4  g0785(.a(n900), .b(n750), .c(n844), .d(in32), .O(n901));
  nand3  g0786(.a(n901), .b(n897), .c(n288), .O(n902));
  nand3  g0787(.a(n902), .b(n509), .c(in26), .O(n903));
  xnor2a g0788(.a(n903), .b(n613), .O(n904));
  nand3  g0789(.a(n904), .b(n440), .c(in36), .O(n905));
  xor2a  g0790(.a(n905), .b(n817), .O(n906));
  nand4  g0791(.a(n906), .b(n896), .c(n895), .d(n787), .O(n907));
  nand3  g0792(.a(n896), .b(n895), .c(n787), .O(n908));
  not    g0793(.a(n906), .O(n909));
  nand2  g0794(.a(n909), .b(n908), .O(n910));
  or2    g0795(.a(n723), .b(in19), .O(n911));
  not    g0796(.a(n911), .O(n912));
  nand3  g0797(.a(n912), .b(n910), .c(n907), .O(n913));
  nand3  g0798(.a(n900), .b(n699), .c(n370), .O(n914));
  nand2  g0799(.a(n914), .b(n358), .O(n915));
  nand3  g0800(.a(n915), .b(n737), .c(n242), .O(n916));
  xor2a  g0801(.a(n643), .b(n557), .O(n917));
  xor2a  g0802(.a(n917), .b(n916), .O(n918));
  nand2  g0803(.a(n918), .b(n639), .O(n919));
  and2   g0804(.a(n919), .b(n201), .O(n920));
  xor2a  g0805(.a(n791), .b(n585), .O(n921));
  nor2   g0806(.a(n921), .b(n185), .O(n922));
  nand4  g0807(.a(n922), .b(n920), .c(n913), .d(n786), .O(n923));
  xor2a  g0808(.a(n745), .b(n168), .O(n924));
  xor2a  g0809(.a(n924), .b(n923), .O(n925));
  or2    g0810(.a(n655), .b(n169), .O(n926));
  nor2   g0811(.a(n926), .b(n925), .O(n927));
  not    g0812(.a(n860), .O(n928));
  not    g0813(.a(n771), .O(n929));
  not    g0814(.a(n601), .O(n930));
  not    g0815(.a(n570), .O(n931));
  nand3  g0816(.a(n874), .b(n361), .c(n793), .O(n932));
  nand2  g0817(.a(n875), .b(n276), .O(n933));
  not    g0818(.a(n760), .O(n934));
  or2    g0819(.a(n934), .b(in72), .O(n935));
  not    g0820(.a(n935), .O(n936));
  nand3  g0821(.a(n936), .b(n933), .c(n932), .O(n937));
  nand2  g0822(.a(n937), .b(n693), .O(n938));
  not    g0823(.a(n814), .O(n939));
  or2    g0824(.a(n939), .b(n424), .O(n940));
  not    g0825(.a(n940), .O(n941));
  nand2  g0826(.a(n941), .b(n938), .O(n942));
  xor2a  g0827(.a(n942), .b(n931), .O(n943));
  xor2a  g0828(.a(n519), .b(n345), .O(n944));
  nand3  g0829(.a(n944), .b(n943), .c(n484), .O(n945));
  nand2  g0830(.a(n943), .b(n484), .O(n946));
  not    g0831(.a(n944), .O(n947));
  nand2  g0832(.a(n947), .b(n946), .O(n948));
  nand2  g0833(.a(n904), .b(n861), .O(n949));
  and2   g0834(.a(n949), .b(in6), .O(n950));
  nand3  g0835(.a(n950), .b(n948), .c(n945), .O(n951));
  nand3  g0836(.a(n951), .b(n930), .c(n929), .O(n952));
  nand2  g0837(.a(n952), .b(n928), .O(n953));
  nand4  g0838(.a(n951), .b(n860), .c(n930), .d(n929), .O(n954));
  and2   g0839(.a(n904), .b(n155), .O(n955));
  nand3  g0840(.a(n955), .b(n954), .c(n953), .O(n956));
  or2    g0841(.a(n956), .b(n927), .O(n957));
  not    g0842(.a(n186), .O(n958));
  or2    g0843(.a(n721), .b(n958), .O(n959));
  not    g0844(.a(n959), .O(n960));
  nand2  g0845(.a(n960), .b(n957), .O(n961));
  not    g0846(.a(n961), .O(n962));
  not    g0847(.a(n522), .O(n963));
  nand3  g0848(.a(n905), .b(n613), .c(n291), .O(n964));
  nand2  g0849(.a(n964), .b(n805), .O(n965));
  xnor2a g0850(.a(n965), .b(n919), .O(n966));
  nand3  g0851(.a(n966), .b(n594), .c(n798), .O(n967));
  not    g0852(.a(n509), .O(n968));
  not    g0853(.a(n592), .O(n969));
  not    g0854(.a(n561), .O(n970));
  xor2a  g0855(.a(n745), .b(in20), .O(n971));
  not    g0856(.a(n971), .O(n972));
  xor2a  g0857(.a(n972), .b(n919), .O(n973));
  not    g0858(.a(in2), .O(n974));
  and2   g0859(.a(n769), .b(n974), .O(n975));
  nand4  g0860(.a(n975), .b(n973), .c(n663), .d(in23), .O(n976));
  nand2  g0861(.a(n976), .b(n970), .O(n977));
  nand4  g0862(.a(n977), .b(n969), .c(n968), .d(n761), .O(n978));
  xor2a  g0863(.a(n607), .b(n313), .O(n979));
  xor2a  g0864(.a(n979), .b(n978), .O(n980));
  nand2  g0865(.a(n980), .b(n739), .O(n981));
  nand2  g0866(.a(n981), .b(n967), .O(n982));
  xor2a  g0867(.a(n592), .b(n465), .O(n983));
  xnor2a g0868(.a(n983), .b(n982), .O(n984));
  not    g0869(.a(n984), .O(n985));
  not    g0870(.a(n518), .O(n986));
  not    g0871(.a(n857), .O(n987));
  nand3  g0872(.a(n949), .b(n987), .c(n986), .O(n988));
  xor2a  g0873(.a(n988), .b(n640), .O(n989));
  nand4  g0874(.a(n989), .b(n985), .c(n714), .d(n709), .O(n990));
  nand3  g0875(.a(n985), .b(n714), .c(n709), .O(n991));
  not    g0876(.a(n989), .O(n992));
  nand2  g0877(.a(n992), .b(n991), .O(n993));
  or2    g0878(.a(n805), .b(n172), .O(n994));
  not    g0879(.a(n994), .O(n995));
  nand3  g0880(.a(n995), .b(n993), .c(n990), .O(n996));
  or2    g0881(.a(n829), .b(n684), .O(n997));
  not    g0882(.a(n997), .O(n998));
  not    g0883(.a(n280), .O(n999));
  and2   g0884(.a(n721), .b(n999), .O(n1000));
  nand4  g0885(.a(n1000), .b(n998), .c(n996), .d(n799), .O(n1001));
  and2   g0886(.a(n769), .b(n117), .O(n1002));
  and2   g0887(.a(n1002), .b(n1001), .O(n1003));
  not    g0888(.a(n1003), .O(n1004));
  not    g0889(.a(n675), .O(n1005));
  not    g0890(.a(n745), .O(n1006));
  nand3  g0891(.a(n1002), .b(n1001), .c(n1006), .O(n1007));
  not    g0892(.a(n1007), .O(n1008));
  not    g0893(.a(n749), .O(n1009));
  and2   g0894(.a(n1009), .b(n425), .O(n1010));
  and2   g0895(.a(n631), .b(n166), .O(n1011));
  nand3  g0896(.a(n1011), .b(n1010), .c(n1008), .O(n1012));
  nand2  g0897(.a(n1012), .b(n1005), .O(n1013));
  xor2a  g0898(.a(n802), .b(n155), .O(n1014));
  not    g0899(.a(n1014), .O(n1015));
  xor2a  g0900(.a(n1015), .b(n1013), .O(n1016));
  not    g0901(.a(n520), .O(n1017));
  nand2  g0902(.a(n1014), .b(n1013), .O(n1018));
  nand3  g0903(.a(n1015), .b(n1012), .c(n1005), .O(n1019));
  or2    g0904(.a(n519), .b(n556), .O(n1020));
  not    g0905(.a(n1020), .O(n1021));
  nand3  g0906(.a(n1021), .b(n1019), .c(n1018), .O(n1022));
  nand2  g0907(.a(n1022), .b(n853), .O(n1023));
  not    g0908(.a(n652), .O(n1024));
  not    g0909(.a(n650), .O(n1025));
  nand3  g0910(.a(n967), .b(n1025), .c(in104), .O(n1026));
  not    g0911(.a(n590), .O(n1027));
  or2    g0912(.a(n1026), .b(n701), .O(n1028));
  nand3  g0913(.a(n1028), .b(n1027), .c(n236), .O(n1029));
  xor2a  g0914(.a(n1029), .b(n778), .O(n1030));
  nand3  g0915(.a(n1030), .b(n1026), .c(n1024), .O(n1031));
  xor2a  g0916(.a(n796), .b(in59), .O(n1032));
  xor2a  g0917(.a(n1032), .b(n1031), .O(n1033));
  xnor2a g0918(.a(n154), .b(n127), .O(n1034));
  xor2a  g0919(.a(n874), .b(n1034), .O(n1035));
  nand3  g0920(.a(n1035), .b(n1033), .c(n537), .O(n1036));
  nand2  g0921(.a(n1033), .b(n537), .O(n1037));
  not    g0922(.a(n1035), .O(n1038));
  nand2  g0923(.a(n1038), .b(n1037), .O(n1039));
  nand3  g0924(.a(n1039), .b(n1036), .c(n400), .O(n1040));
  not    g0925(.a(n1040), .O(n1041));
  nand4  g0926(.a(n1041), .b(n1023), .c(n915), .d(n999), .O(n1042));
  nand3  g0927(.a(n1041), .b(n1023), .c(n999), .O(n1043));
  nand3  g0928(.a(n1043), .b(n914), .c(n358), .O(n1044));
  and2   g0929(.a(n1007), .b(in78), .O(n1045));
  nand4  g0930(.a(n1045), .b(n1044), .c(n1042), .d(n1012), .O(n1046));
  xor2a  g0931(.a(n851), .b(in59), .O(n1047));
  xor2a  g0932(.a(n1047), .b(n956), .O(n1048));
  nand3  g0933(.a(n977), .b(n969), .c(n443), .O(n1049));
  not    g0934(.a(n1049), .O(n1050));
  nand2  g0935(.a(n1050), .b(n1048), .O(n1051));
  xor2a  g0936(.a(n1033), .b(n551), .O(n1052));
  xor2a  g0937(.a(n1052), .b(n1051), .O(n1053));
  or2    g0938(.a(n1007), .b(n764), .O(n1054));
  not    g0939(.a(n1054), .O(n1055));
  nand2  g0940(.a(n1055), .b(n1053), .O(n1056));
  xor2a  g0941(.a(n1056), .b(n1046), .O(n1057));
  not    g0942(.a(n851), .O(n1058));
  not    g0943(.a(n1001), .O(n1059));
  not    g0944(.a(n856), .O(n1060));
  nand2  g0945(.a(n975), .b(n973), .O(n1061));
  not    g0946(.a(n1061), .O(n1062));
  nand4  g0947(.a(n1057), .b(n922), .c(n920), .d(n913), .O(n1063));
  nand2  g0948(.a(n1063), .b(n891), .O(n1064));
  nand2  g0949(.a(n1064), .b(n657), .O(n1065));
  xor2a  g0950(.a(n1065), .b(n1062), .O(n1066));
  or2    g0951(.a(n996), .b(in109), .O(n1067));
  not    g0952(.a(n1067), .O(n1068));
  nand2  g0953(.a(n1068), .b(n1066), .O(n1069));
  not    g0954(.a(n551), .O(n1070));
  and2   g0955(.a(n942), .b(n1070), .O(n1071));
  nand3  g0956(.a(n1071), .b(n1069), .c(n1060), .O(n1072));
  nand2  g0957(.a(n1072), .b(n668), .O(n1073));
  or2    g0958(.a(n596), .b(in80), .O(n1074));
  not    g0959(.a(n1074), .O(n1075));
  nand2  g0960(.a(n1075), .b(n1073), .O(n1076));
  xor2a  g0961(.a(n656), .b(n211), .O(n1077));
  nand2  g0962(.a(n1077), .b(n1076), .O(n1078));
  not    g0963(.a(n1077), .O(n1079));
  nand3  g0964(.a(n1079), .b(n1075), .c(n1073), .O(n1080));
  nand3  g0965(.a(n1080), .b(n1078), .c(n706), .O(n1081));
  nand2  g0966(.a(n1081), .b(n564), .O(n1082));
  nand2  g0967(.a(n1082), .b(n1059), .O(n1083));
  xor2a  g0968(.a(n1083), .b(n1058), .O(n1084));
  nand2  g0969(.a(n1084), .b(n757), .O(n1085));
  xor2a  g0970(.a(n1083), .b(n851), .O(n1086));
  nand2  g0971(.a(n1086), .b(n756), .O(n1087));
  or2    g0972(.a(n1013), .b(in19), .O(n1088));
  not    g0973(.a(n1088), .O(n1089));
  nand3  g0974(.a(n1089), .b(n1087), .c(n1085), .O(n1090));
  nand2  g0975(.a(n1090), .b(n1057), .O(n1091));
  nand2  g0976(.a(n1091), .b(n1017), .O(n1092));
  xor2a  g0977(.a(n1092), .b(n1016), .O(n1093));
  and2   g0978(.a(n905), .b(n291), .O(n1094));
  not    g0979(.a(n565), .O(n1095));
  or2    g0980(.a(n988), .b(n852), .O(n1096));
  nand3  g0981(.a(n1096), .b(n728), .c(n1095), .O(n1097));
  not    g0982(.a(n1097), .O(n1098));
  nand3  g0983(.a(n1098), .b(n856), .c(n458), .O(n1099));
  xor2a  g0984(.a(n1099), .b(n590), .O(n1100));
  nor3   g0985(.a(n1100), .b(n1094), .c(n493), .O(n1101));
  xnor2a g0986(.a(n908), .b(in88), .O(n1102));
  xor2a  g0987(.a(n1102), .b(n1101), .O(n1103));
  and2   g0988(.a(n998), .b(n996), .O(n1104));
  nand4  g0989(.a(n1055), .b(n1053), .c(n1104), .d(n799), .O(n1105));
  and2   g0990(.a(n1105), .b(n1103), .O(n1106));
  xnor2a g0991(.a(n1106), .b(n735), .O(n1107));
  or2    g0992(.a(n1043), .b(n432), .O(n1108));
  or2    g0993(.a(n1108), .b(n1107), .O(n1109));
  or2    g0994(.a(n1109), .b(in4), .O(n1110));
  not    g0995(.a(n1110), .O(n1111));
  nand4  g0996(.a(n1111), .b(n1093), .c(n1004), .d(n963), .O(n1112));
  xor2a  g0997(.a(n1112), .b(n706), .O(n1113));
  xor2a  g0998(.a(n1113), .b(n757), .O(n1114));
  xor2a  g0999(.a(n952), .b(n311), .O(n1115));
  xor2a  g1000(.a(n1115), .b(n1114), .O(n1116));
  nand2  g1001(.a(n1116), .b(n538), .O(n1117));
  not    g1002(.a(n538), .O(n1118));
  xor2a  g1003(.a(n1113), .b(n756), .O(n1119));
  xor2a  g1004(.a(n1115), .b(n1119), .O(n1120));
  nand2  g1005(.a(n1120), .b(n1118), .O(n1121));
  not    g1006(.a(n741), .O(n1122));
  not    g1007(.a(n370), .O(n1123));
  not    g1008(.a(n996), .O(n1124));
  not    g1009(.a(n949), .O(n1125));
  or2    g1010(.a(n1125), .b(n518), .O(n1126));
  nand2  g1011(.a(n779), .b(n777), .O(n1127));
  not    g1012(.a(n605), .O(n1128));
  not    g1013(.a(n403), .O(n1129));
  nand3  g1014(.a(n1103), .b(n966), .c(n1129), .O(n1130));
  nand4  g1015(.a(n1130), .b(n914), .c(n724), .d(n152), .O(n1131));
  xor2a  g1016(.a(n594), .b(in35), .O(n1132));
  xor2a  g1017(.a(n1132), .b(n1131), .O(n1133));
  nand4  g1018(.a(n1133), .b(n1128), .c(n1127), .d(n214), .O(n1134));
  or2    g1019(.a(n1134), .b(n736), .O(n1135));
  not    g1020(.a(n1135), .O(n1136));
  or2    g1021(.a(n1136), .b(n1126), .O(n1137));
  and2   g1022(.a(n1137), .b(n624), .O(n1138));
  xnor2a g1023(.a(n923), .b(in41), .O(n1139));
  xor2a  g1024(.a(n1139), .b(n1138), .O(n1140));
  nand3  g1025(.a(n1140), .b(n1124), .c(n1122), .O(n1141));
  nand3  g1026(.a(n1141), .b(n655), .c(n775), .O(n1142));
  not    g1027(.a(n653), .O(n1143));
  not    g1028(.a(n237), .O(n1144));
  xor2a  g1029(.a(n894), .b(n891), .O(n1145));
  not    g1030(.a(n927), .O(n1146));
  not    g1031(.a(n859), .O(n1147));
  nand4  g1032(.a(n961), .b(n748), .c(n747), .d(in1), .O(n1148));
  nand3  g1033(.a(n1148), .b(n1147), .c(n261), .O(n1149));
  nand3  g1034(.a(n1149), .b(n1146), .c(n666), .O(n1150));
  nand2  g1035(.a(n1150), .b(n921), .O(n1151));
  and2   g1036(.a(n1100), .b(n171), .O(n1152));
  and2   g1037(.a(n1152), .b(n1151), .O(n1153));
  or2    g1038(.a(n919), .b(n164), .O(n1154));
  not    g1039(.a(n1154), .O(n1155));
  nand4  g1040(.a(n1155), .b(n1153), .c(n1145), .d(n1144), .O(n1156));
  nand3  g1041(.a(n1156), .b(n880), .c(n879), .O(n1157));
  xor2a  g1042(.a(n1126), .b(n125), .O(n1158));
  xor2a  g1043(.a(n1158), .b(n1157), .O(n1159));
  or2    g1044(.a(n1159), .b(n1143), .O(n1160));
  nand3  g1045(.a(n1160), .b(n1059), .c(n262), .O(n1161));
  not    g1046(.a(n883), .O(n1162));
  or2    g1047(.a(n1162), .b(n496), .O(n1163));
  not    g1048(.a(n1163), .O(n1164));
  nand4  g1049(.a(n1164), .b(n1161), .c(n1142), .d(n1123), .O(n1165));
  and2   g1050(.a(n976), .b(in51), .O(n1166));
  nand3  g1051(.a(n1166), .b(n1165), .c(n1122), .O(n1167));
  xor2a  g1052(.a(n1167), .b(n879), .O(n1168));
  and2   g1053(.a(n1151), .b(n372), .O(n1169));
  and2   g1054(.a(n1001), .b(n215), .O(n1170));
  nand4  g1055(.a(n1170), .b(n1169), .c(n1168), .d(n568), .O(n1171));
  not    g1056(.a(n1171), .O(n1172));
  not    g1057(.a(in55), .O(n1173));
  nor2   g1058(.a(n984), .b(n706), .O(n1174));
  not    g1059(.a(n791), .O(n1175));
  xor2a  g1060(.a(n752), .b(in56), .O(n1176));
  xor2a  g1061(.a(n1176), .b(n1040), .O(n1177));
  xor2a  g1062(.a(n1177), .b(n291), .O(n1178));
  nand2  g1063(.a(n1178), .b(n1175), .O(n1179));
  nand3  g1064(.a(n1179), .b(n1003), .c(in10), .O(n1180));
  xor2a  g1065(.a(n411), .b(n556), .O(n1181));
  xor2a  g1066(.a(n1181), .b(n1180), .O(n1182));
  xor2a  g1067(.a(n1182), .b(n1098), .O(n1183));
  xor2a  g1068(.a(n903), .b(in61), .O(n1184));
  xor2a  g1069(.a(n1184), .b(n1183), .O(n1185));
  nand4  g1070(.a(n1185), .b(n964), .c(n805), .d(n192), .O(n1186));
  nand3  g1071(.a(n1186), .b(n976), .c(n970), .O(n1187));
  nand3  g1072(.a(n1187), .b(n668), .c(n1009), .O(n1188));
  nand2  g1073(.a(n1188), .b(n814), .O(n1189));
  xor2a  g1074(.a(n1189), .b(n1174), .O(n1190));
  nand3  g1075(.a(n889), .b(n866), .c(in7), .O(n1191));
  or2    g1076(.a(n982), .b(n195), .O(n1192));
  not    g1077(.a(n1192), .O(n1193));
  nand4  g1078(.a(n1193), .b(n1191), .c(n916), .d(n557), .O(n1194));
  xor2a  g1079(.a(n991), .b(n248), .O(n1195));
  xor2a  g1080(.a(n1195), .b(n1194), .O(n1196));
  xor2a  g1081(.a(n1196), .b(in51), .O(n1197));
  xor2a  g1082(.a(n1197), .b(n1190), .O(n1198));
  nand4  g1083(.a(n1198), .b(n802), .c(n733), .d(n485), .O(n1199));
  nand3  g1084(.a(n1199), .b(n1030), .c(n186), .O(n1200));
  or2    g1085(.a(n1200), .b(n1173), .O(n1201));
  not    g1086(.a(n1201), .O(n1202));
  nand4  g1087(.a(n1202), .b(n1172), .c(n1121), .d(n1117), .O(n1203));
  and2   g1088(.a(n1187), .b(n187), .O(n1204));
  nand2  g1089(.a(n1204), .b(n1203), .O(n1205));
  xor2a  g1090(.a(n1205), .b(n1113), .O(n1206));
  xor2a  g1091(.a(n1109), .b(in60), .O(n1207));
  xor2a  g1092(.a(n1207), .b(n1206), .O(n1208));
  nor2   g1093(.a(n725), .b(n156), .O(n1209));
  or2    g1094(.a(n1185), .b(n496), .O(n1210));
  not    g1095(.a(n1210), .O(n1211));
  nand4  g1096(.a(n1211), .b(n1209), .c(n1208), .d(n962), .O(n1212));
  not    g1097(.a(n1161), .O(n1213));
  not    g1098(.a(n1188), .O(n1214));
  nor4   g1099(.a(n1194), .b(n1108), .c(n1107), .d(n303), .O(n1215));
  or2    g1100(.a(n1215), .b(n1214), .O(n1216));
  and2   g1101(.a(n1030), .b(n1026), .O(n1217));
  xor2a  g1102(.a(n1217), .b(n190), .O(n1218));
  xor2a  g1103(.a(n1218), .b(n1216), .O(n1219));
  or2    g1104(.a(n1219), .b(n482), .O(n1220));
  xnor2a g1105(.a(n1189), .b(in18), .O(n1221));
  xor2a  g1106(.a(n1221), .b(n1220), .O(n1222));
  nand4  g1107(.a(n1222), .b(n1213), .c(n298), .d(in64), .O(n1223));
  xor2a  g1108(.a(n1097), .b(n389), .O(n1224));
  xor2a  g1109(.a(n1224), .b(n1223), .O(n1225));
  nand4  g1110(.a(n1225), .b(n1044), .c(n1042), .d(in56), .O(n1226));
  and2   g1111(.a(n1226), .b(n239), .O(n1227));
  not    g1112(.a(n908), .O(n1228));
  xor2a  g1113(.a(n1200), .b(n1190), .O(n1229));
  xor2a  g1114(.a(n881), .b(n308), .O(n1230));
  nand2  g1115(.a(n1230), .b(n1229), .O(n1231));
  not    g1116(.a(n1190), .O(n1232));
  xor2a  g1117(.a(n1200), .b(n1232), .O(n1233));
  not    g1118(.a(n1230), .O(n1234));
  nand2  g1119(.a(n1234), .b(n1233), .O(n1235));
  nand3  g1120(.a(n1235), .b(n1231), .c(n988), .O(n1236));
  nand3  g1121(.a(n1236), .b(n925), .c(n178), .O(n1237));
  xor2a  g1122(.a(n1237), .b(n1134), .O(n1238));
  nand2  g1123(.a(n1238), .b(n787), .O(n1239));
  nand2  g1124(.a(n1239), .b(n1006), .O(n1240));
  not    g1125(.a(n250), .O(n1241));
  or2    g1126(.a(n1066), .b(n1241), .O(n1242));
  not    g1127(.a(n1242), .O(n1243));
  nand4  g1128(.a(n1243), .b(n1240), .c(n1029), .d(n495), .O(n1244));
  nand2  g1129(.a(n1244), .b(n626), .O(n1245));
  nand2  g1130(.a(n1245), .b(n1012), .O(n1246));
  not    g1131(.a(n1012), .O(n1247));
  nand3  g1132(.a(n1244), .b(n1247), .c(n626), .O(n1248));
  nand3  g1133(.a(n1248), .b(n1246), .c(n851), .O(n1249));
  xnor2a g1134(.a(n1249), .b(n1046), .O(n1250));
  nand3  g1135(.a(n1250), .b(n1007), .c(n219), .O(n1251));
  nand2  g1136(.a(n1251), .b(n1165), .O(n1252));
  xor2a  g1137(.a(n1252), .b(n1228), .O(n1253));
  nand2  g1138(.a(n1253), .b(n791), .O(n1254));
  xor2a  g1139(.a(n1252), .b(n908), .O(n1255));
  nand2  g1140(.a(n1255), .b(n1175), .O(n1256));
  nand3  g1141(.a(n1256), .b(n1254), .c(n150), .O(n1257));
  not    g1142(.a(n1257), .O(n1258));
  nand3  g1143(.a(n1258), .b(n1227), .c(n1212), .O(n1259));
  not    g1144(.a(n431), .O(n1260));
  and2   g1145(.a(n1189), .b(n1260), .O(n1261));
  nand2  g1146(.a(n1261), .b(n1259), .O(n1262));
  nand2  g1147(.a(n1262), .b(n890), .O(out1));
endmodule


