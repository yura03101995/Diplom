module mux_9 ( ctrl0, ctrl1, ctrl2, ctrl3, ctrl4, ctrl5, ctrl6, ctrl7, ctrl8, in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, in64, in65, in66, in67, in68, in69, in70, in71, in72, in73, in74, in75, in76, in77, in78, in79, in80, in81, in82, in83, in84, in85, in86, in87, in88, in89, in90, in91, in92, in93, in94, in95, in96, in97, in98, in99, in100, in101, in102, in103, in104, in105, in106, in107, in108, in109, in110, in111, in112, in113, in114, in115, in116, in117, in118, in119, in120, in121, in122, in123, in124, in125, in126, in127, in128, in129, in130, in131, in132, in133, in134, in135, in136, in137, in138, in139, in140, in141, in142, in143, in144, in145, in146, in147, in148, in149, in150, in151, in152, in153, in154, in155, in156, in157, in158, in159, in160, in161, in162, in163, in164, in165, in166, in167, in168, in169, in170, in171, in172, in173, in174, in175, in176, in177, in178, in179, in180, in181, in182, in183, in184, in185, in186, in187, in188, in189, in190, in191, in192, in193, in194, in195, in196, in197, in198, in199, in200, in201, in202, in203, in204, in205, in206, in207, in208, in209, in210, in211, in212, in213, in214, in215, in216, in217, in218, in219, in220, in221, in222, in223, in224, in225, in226, in227, in228, in229, in230, in231, in232, in233, in234, in235, in236, in237, in238, in239, in240, in241, in242, in243, in244, in245, in246, in247, in248, in249, in250, in251, in252, in253, in254, in255, in256, in257, in258, in259, in260, in261, in262, in263, in264, in265, in266, in267, in268, in269, in270, in271, in272, in273, in274, in275, in276, in277, in278, in279, in280, in281, in282, in283, in284, in285, in286, in287, in288, in289, in290, in291, in292, in293, in294, in295, in296, in297, in298, in299, in300, in301, in302, in303, in304, in305, in306, in307, in308, in309, in310, in311, in312, in313, in314, in315, in316, in317, in318, in319, in320, in321, in322, in323, in324, in325, in326, in327, in328, in329, in330, in331, in332, in333, in334, in335, in336, in337, in338, in339, in340, in341, in342, in343, in344, in345, in346, in347, in348, in349, in350, in351, in352, in353, in354, in355, in356, in357, in358, in359, in360, in361, in362, in363, in364, in365, in366, in367, in368, in369, in370, in371, in372, in373, in374, in375, in376, in377, in378, in379, in380, in381, in382, in383, in384, in385, in386, in387, in388, in389, in390, in391, in392, in393, in394, in395, in396, in397, in398, in399, in400, in401, in402, in403, in404, in405, in406, in407, in408, in409, in410, in411, in412, in413, in414, in415, in416, in417, in418, in419, in420, in421, in422, in423, in424, in425, in426, in427, in428, in429, in430, in431, in432, in433, in434, in435, in436, in437, in438, in439, in440, in441, in442, in443, in444, in445, in446, in447, in448, in449, in450, in451, in452, in453, in454, in455, in456, in457, in458, in459, in460, in461, in462, in463, in464, in465, in466, in467, in468, in469, in470, in471, in472, in473, in474, in475, in476, in477, in478, in479, in480, in481, in482, in483, in484, in485, in486, in487, in488, in489, in490, in491, in492, in493, in494, in495, in496, in497, in498, in499, in500, in501, in502, in503, in504, in505, in506, in507, in508, in509, in510, in511, out);
input ctrl0, ctrl1, ctrl2, ctrl3, ctrl4, ctrl5, ctrl6, ctrl7, ctrl8, in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, in64, in65, in66, in67, in68, in69, in70, in71, in72, in73, in74, in75, in76, in77, in78, in79, in80, in81, in82, in83, in84, in85, in86, in87, in88, in89, in90, in91, in92, in93, in94, in95, in96, in97, in98, in99, in100, in101, in102, in103, in104, in105, in106, in107, in108, in109, in110, in111, in112, in113, in114, in115, in116, in117, in118, in119, in120, in121, in122, in123, in124, in125, in126, in127, in128, in129, in130, in131, in132, in133, in134, in135, in136, in137, in138, in139, in140, in141, in142, in143, in144, in145, in146, in147, in148, in149, in150, in151, in152, in153, in154, in155, in156, in157, in158, in159, in160, in161, in162, in163, in164, in165, in166, in167, in168, in169, in170, in171, in172, in173, in174, in175, in176, in177, in178, in179, in180, in181, in182, in183, in184, in185, in186, in187, in188, in189, in190, in191, in192, in193, in194, in195, in196, in197, in198, in199, in200, in201, in202, in203, in204, in205, in206, in207, in208, in209, in210, in211, in212, in213, in214, in215, in216, in217, in218, in219, in220, in221, in222, in223, in224, in225, in226, in227, in228, in229, in230, in231, in232, in233, in234, in235, in236, in237, in238, in239, in240, in241, in242, in243, in244, in245, in246, in247, in248, in249, in250, in251, in252, in253, in254, in255, in256, in257, in258, in259, in260, in261, in262, in263, in264, in265, in266, in267, in268, in269, in270, in271, in272, in273, in274, in275, in276, in277, in278, in279, in280, in281, in282, in283, in284, in285, in286, in287, in288, in289, in290, in291, in292, in293, in294, in295, in296, in297, in298, in299, in300, in301, in302, in303, in304, in305, in306, in307, in308, in309, in310, in311, in312, in313, in314, in315, in316, in317, in318, in319, in320, in321, in322, in323, in324, in325, in326, in327, in328, in329, in330, in331, in332, in333, in334, in335, in336, in337, in338, in339, in340, in341, in342, in343, in344, in345, in346, in347, in348, in349, in350, in351, in352, in353, in354, in355, in356, in357, in358, in359, in360, in361, in362, in363, in364, in365, in366, in367, in368, in369, in370, in371, in372, in373, in374, in375, in376, in377, in378, in379, in380, in381, in382, in383, in384, in385, in386, in387, in388, in389, in390, in391, in392, in393, in394, in395, in396, in397, in398, in399, in400, in401, in402, in403, in404, in405, in406, in407, in408, in409, in410, in411, in412, in413, in414, in415, in416, in417, in418, in419, in420, in421, in422, in423, in424, in425, in426, in427, in428, in429, in430, in431, in432, in433, in434, in435, in436, in437, in438, in439, in440, in441, in442, in443, in444, in445, in446, in447, in448, in449, in450, in451, in452, in453, in454, in455, in456, in457, in458, in459, in460, in461, in462, in463, in464, in465, in466, in467, in468, in469, in470, in471, in472, in473, in474, in475, in476, in477, in478, in479, in480, in481, in482, in483, in484, in485, in486, in487, in488, in489, in490, in491, in492, in493, in494, in495, in496, in497, in498, in499, in500, in501, in502, in503, in504, in505, in506, in507, in508, in509, in510, in511;
output out;
assign out = ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in1 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in2 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in3 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in4 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in5 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in6 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in7 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in8 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in9 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in10 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in11 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in12 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in13 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in14 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in15 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in16 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in17 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in18 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in19 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in20 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in21 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in22 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in23 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in24 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in25 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in26 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in27 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in28 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in29 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in30 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in31 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in32 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in33 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in34 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in35 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in36 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in37 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in38 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in39 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in40 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in41 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in42 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in43 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in44 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in45 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in46 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in47 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in48 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in49 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in50 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in51 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in52 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in53 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in54 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in55 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in56 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in57 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in58 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in59 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in60 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in61 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in62 : 
             ( ~ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in63 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in64 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in65 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in66 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in67 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in68 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in69 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in70 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in71 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in72 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in73 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in74 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in75 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in76 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in77 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in78 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in79 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in80 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in81 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in82 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in83 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in84 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in85 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in86 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in87 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in88 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in89 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in90 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in91 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in92 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in93 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in94 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in95 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in96 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in97 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in98 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in99 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in100 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in101 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in102 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in103 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in104 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in105 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in106 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in107 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in108 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in109 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in110 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in111 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in112 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in113 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in114 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in115 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in116 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in117 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in118 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in119 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in120 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in121 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in122 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in123 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in124 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in125 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in126 : 
             ( ~ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in127 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in128 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in129 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in130 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in131 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in132 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in133 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in134 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in135 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in136 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in137 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in138 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in139 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in140 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in141 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in142 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in143 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in144 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in145 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in146 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in147 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in148 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in149 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in150 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in151 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in152 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in153 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in154 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in155 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in156 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in157 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in158 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in159 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in160 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in161 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in162 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in163 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in164 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in165 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in166 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in167 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in168 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in169 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in170 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in171 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in172 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in173 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in174 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in175 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in176 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in177 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in178 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in179 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in180 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in181 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in182 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in183 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in184 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in185 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in186 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in187 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in188 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in189 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in190 : 
             ( ~ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in191 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in192 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in193 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in194 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in195 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in196 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in197 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in198 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in199 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in200 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in201 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in202 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in203 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in204 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in205 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in206 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in207 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in208 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in209 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in210 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in211 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in212 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in213 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in214 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in215 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in216 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in217 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in218 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in219 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in220 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in221 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in222 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in223 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in224 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in225 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in226 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in227 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in228 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in229 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in230 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in231 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in232 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in233 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in234 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in235 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in236 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in237 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in238 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in239 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in240 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in241 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in242 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in243 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in244 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in245 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in246 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in247 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in248 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in249 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in250 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in251 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in252 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in253 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in254 : 
             ( ~ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in255 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in256 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in257 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in258 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in259 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in260 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in261 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in262 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in263 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in264 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in265 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in266 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in267 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in268 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in269 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in270 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in271 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in272 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in273 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in274 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in275 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in276 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in277 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in278 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in279 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in280 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in281 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in282 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in283 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in284 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in285 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in286 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in287 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in288 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in289 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in290 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in291 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in292 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in293 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in294 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in295 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in296 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in297 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in298 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in299 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in300 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in301 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in302 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in303 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in304 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in305 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in306 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in307 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in308 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in309 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in310 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in311 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in312 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in313 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in314 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in315 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in316 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in317 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in318 : 
             ( ctrl0 & ~ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in319 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in320 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in321 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in322 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in323 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in324 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in325 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in326 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in327 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in328 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in329 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in330 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in331 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in332 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in333 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in334 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in335 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in336 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in337 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in338 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in339 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in340 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in341 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in342 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in343 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in344 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in345 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in346 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in347 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in348 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in349 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in350 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in351 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in352 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in353 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in354 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in355 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in356 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in357 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in358 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in359 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in360 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in361 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in362 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in363 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in364 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in365 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in366 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in367 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in368 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in369 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in370 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in371 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in372 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in373 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in374 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in375 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in376 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in377 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in378 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in379 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in380 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in381 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in382 : 
             ( ctrl0 & ~ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in383 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in384 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in385 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in386 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in387 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in388 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in389 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in390 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in391 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in392 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in393 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in394 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in395 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in396 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in397 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in398 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in399 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in400 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in401 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in402 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in403 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in404 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in405 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in406 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in407 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in408 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in409 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in410 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in411 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in412 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in413 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in414 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in415 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in416 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in417 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in418 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in419 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in420 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in421 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in422 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in423 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in424 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in425 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in426 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in427 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in428 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in429 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in430 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in431 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in432 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in433 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in434 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in435 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in436 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in437 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in438 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in439 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in440 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in441 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in442 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in443 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in444 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in445 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in446 : 
             ( ctrl0 & ctrl1 & ~ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in447 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in448 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in449 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in450 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in451 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in452 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in453 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in454 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in455 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in456 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in457 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in458 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in459 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in460 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in461 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in462 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in463 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in464 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in465 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in466 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in467 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in468 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in469 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in470 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in471 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in472 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in473 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in474 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in475 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in476 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in477 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in478 : 
             ( ctrl0 & ctrl1 & ctrl2 & ~ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in479 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in480 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in481 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in482 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in483 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in484 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in485 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in486 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in487 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in488 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in489 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in490 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in491 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in492 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in493 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in494 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ~ctrl4 & ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in495 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in496 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in497 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in498 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in499 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in500 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in501 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in502 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ~ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in503 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ~ctrl8  ) ? in504 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ~ctrl7 & ctrl8  ) ? in505 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ~ctrl8  ) ? in506 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ~ctrl6 & ctrl7 & ctrl8  ) ? in507 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ~ctrl8  ) ? in508 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ~ctrl7 & ctrl8  ) ? in509 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7 & ~ctrl8  ) ? in510 : 
             ( ctrl0 & ctrl1 & ctrl2 & ctrl3 & ctrl4 & ctrl5 & ctrl6 & ctrl7 & ctrl8  ) ? in511 : 
             in0;
endmodule
